module background_data(input [18:0] read_address,
								output logic [3:0] value
								);

	assign value = data[read_address];
								
parameter bit [0:307199][2:0] data = {
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h7,
3'h3,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h3,
3'h7,
3'h5,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h7,
3'h7,
3'h7,
3'h3,
3'h2,
3'h2,
3'h3,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h3,
3'h7,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h7,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h7,
3'h7,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h7,
3'h7,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h7,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h5,
3'h7,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h3,
3'h7,
3'h5,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h7,
3'h3,
3'h2,
3'h2,
3'h3,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h3,
3'h7,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h7,
3'h7,
3'h3,
3'h2,
3'h2,
3'h3,
3'h2,
3'h2,
3'h3,
3'h2,
3'h2,
3'h3,
3'h7,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h7,
3'h3,
3'h2,
3'h3,
3'h3,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h3,
3'h7,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h7,
3'h7,
3'h7,
3'h7,
3'h3,
3'h3,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h7,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h7,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h3,
3'h7,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h7,
3'h7,
3'h3,
3'h7,
3'h3,
3'h3,
3'h3,
3'h2,
3'h2,
3'h2,
3'h2,
3'h3,
3'h2,
3'h2,
3'h2,
3'h2,
3'h3,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h7,
3'h7,
3'h3,
3'h3,
3'h7,
3'h7,
3'h7,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h7,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h3,
3'h3,
3'h7,
3'h7,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h7,
3'h7,
3'h7,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h2,
3'h2,
3'h2,
3'h2,
3'h3,
3'h2,
3'h2,
3'h2,
3'h2,
3'h3,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h7,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h3,
3'h5,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h7,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h3,
3'h7,
3'h5,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h7,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h2,
3'h2,
3'h2,
3'h2,
3'h3,
3'h2,
3'h2,
3'h2,
3'h3,
3'h7,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h7,
3'h7,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h7,
3'h7,
3'h7,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h7,
3'h2,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h3,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h5,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h7,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h2,
3'h2,
3'h2,
3'h3,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h7,
3'h3,
3'h3,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h3,
3'h2,
3'h2,
3'h3,
3'h5,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h5,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h3,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h3,
3'h2,
3'h3,
3'h5,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h7,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h7,
3'h3,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h3,
3'h2,
3'h2,
3'h3,
3'h7,
3'h0,
3'h0,
3'h7,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h3,
3'h7,
3'h7,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h7,
3'h7,
3'h3,
3'h2,
3'h3,
3'h3,
3'h2,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h2,
3'h3,
3'h3,
3'h2,
3'h2,
3'h3,
3'h2,
3'h2,
3'h3,
3'h5,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h7,
3'h3,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h3,
3'h2,
3'h2,
3'h7,
3'h0,
3'h0,
3'h7,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h3,
3'h7,
3'h6,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h7,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h3,
3'h5,
3'h5,
3'h5,
3'h7,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h7,
3'h7,
3'h7,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h7,
3'h3,
3'h3,
3'h3,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h3,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h7,
3'h5,
3'h7,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h3,
3'h3,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h3,
3'h7,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h7,
3'h7,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h2,
3'h2,
3'h2,
3'h2,
3'h3,
3'h3,
3'h2,
3'h3,
3'h7,
3'h7,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h5,
3'h7,
3'h7,
3'h3,
3'h7,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h7,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h3,
3'h5,
3'h7,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h7,
3'h7,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h3,
3'h3,
3'h2,
3'h2,
3'h2,
3'h3,
3'h2,
3'h3,
3'h2,
3'h2,
3'h2,
3'h2,
3'h3,
3'h7,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h7,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h2,
3'h2,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h2,
3'h2,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h7,
3'h7,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h5,
3'h7,
3'h3,
3'h3,
3'h3,
3'h3,
3'h7,
3'h7,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h7,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h3,
3'h3,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h3,
3'h2,
3'h2,
3'h2,
3'h2,
3'h3,
3'h7,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h7,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h2,
3'h2,
3'h2,
3'h2,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h2,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h2,
3'h2,
3'h3,
3'h2,
3'h2,
3'h3,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h7,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h3,
3'h7,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h7,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h7,
3'h7,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h5,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h7,
3'h7,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h2,
3'h2,
3'h3,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h3,
3'h3,
3'h3,
3'h2,
3'h2,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h2,
3'h2,
3'h2,
3'h3,
3'h3,
3'h3,
3'h3,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h3,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h7,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h3,
3'h3,
3'h5,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h7,
3'h7,
3'h7,
3'h3,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h3,
3'h7,
3'h7,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h7,
3'h7,
3'h7,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h2,
3'h3,
3'h7,
3'h7,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h5,
3'h3,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h5,
3'h5,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h7,
3'h7,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h2,
3'h3,
3'h3,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h5,
3'h6,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h7,
3'h3,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h5,
3'h5,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h5,
3'h5,
3'h5,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h7,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h7,
3'h7,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h7,
3'h7,
3'h3,
3'h2,
3'h2,
3'h2,
3'h2,
3'h3,
3'h3,
3'h3,
3'h3,
3'h7,
3'h7,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h7,
3'h7,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h2,
3'h3,
3'h2,
3'h2,
3'h3,
3'h2,
3'h2,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h2,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h3,
3'h3,
3'h5,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h3,
3'h2,
3'h3,
3'h3,
3'h7,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h7,
3'h7,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h3,
3'h7,
3'h7,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h7,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h7,
3'h7,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h7,
3'h7,
3'h3,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h7,
3'h7,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h7,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h2,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h2,
3'h3,
3'h3,
3'h5,
3'h3,
3'h2,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h2,
3'h2,
3'h3,
3'h2,
3'h2,
3'h2,
3'h3,
3'h3,
3'h5,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h7,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h2,
3'h2,
3'h2,
3'h2,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h3,
3'h3,
3'h7,
3'h0,
3'h7,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h7,
3'h2,
3'h2,
3'h3,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h3,
3'h7,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h7,
3'h5,
3'h7,
3'h3,
3'h3,
3'h3,
3'h7,
3'h5,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h7,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h7,
3'h7,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h7,
3'h7,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h7,
3'h7,
3'h7,
3'h3,
3'h3,
3'h3,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h7,
3'h7,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h2,
3'h2,
3'h3,
3'h2,
3'h2,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h2,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h7,
3'h5,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h7,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h3,
3'h3,
3'h3,
3'h7,
3'h7,
3'h5,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h5,
3'h7,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h7,
3'h7,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h7,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h7,
3'h7,
3'h7,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h7,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h7,
3'h5,
3'h5,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h7,
3'h7,
3'h7,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h5,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h7,
3'h7,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h2,
3'h3,
3'h3,
3'h3,
3'h2,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h7,
3'h7,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h5,
3'h7,
3'h7,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h5,
3'h2,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h7,
3'h7,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h7,
3'h7,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h2,
3'h7,
3'h7,
3'h7,
3'h7,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h7,
3'h3,
3'h3,
3'h3,
3'h7,
3'h7,
3'h7,
3'h7,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h7,
3'h7,
3'h7,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h7,
3'h7,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h7,
3'h7,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h7,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h3,
3'h3,
3'h3,
3'h3,
3'h2,
3'h3,
3'h3,
3'h7,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h7,
3'h3,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h7,
3'h0,
3'h0,
3'h0,
3'h0,
3'h7,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h7,
3'h2,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h3,
3'h7,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h7,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h7,
3'h7,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h7,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h3,
3'h2,
3'h2,
3'h3,
3'h7,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h7,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h2,
3'h3,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h7,
3'h7,
3'h7,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h7,
3'h3,
3'h2,
3'h3,
3'h3,
3'h2,
3'h2,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h2,
3'h2,
3'h2,
3'h2,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h7,
3'h7,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h7,
3'h7,
3'h7,
3'h3,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h7,
3'h7,
3'h7,
3'h0,
3'h7,
3'h0,
3'h0,
3'h0,
3'h0,
3'h7,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h3,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h7,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h7,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h7,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h2,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h7,
3'h5,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h7,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h2,
3'h2,
3'h2,
3'h3,
3'h3,
3'h3,
3'h2,
3'h3,
3'h3,
3'h7,
3'h7,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h5,
3'h3,
3'h3,
3'h3,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h3,
3'h2,
3'h2,
3'h3,
3'h2,
3'h3,
3'h5,
3'h5,
3'h7,
3'h0,
3'h0,
3'h0,
3'h7,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h3,
3'h3,
3'h7,
3'h0,
3'h7,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h7,
3'h0,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h3,
3'h3,
3'h7,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h5,
3'h7,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h2,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h7,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h7,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h2,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h7,
3'h7,
3'h7,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h5,
3'h3,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h3,
3'h7,
3'h7,
3'h0,
3'h0,
3'h7,
3'h7,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h3,
3'h3,
3'h2,
3'h2,
3'h3,
3'h2,
3'h3,
3'h7,
3'h7,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h5,
3'h5,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h3,
3'h7,
3'h5,
3'h7,
3'h0,
3'h7,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h7,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h7,
3'h7,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h7,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h7,
3'h7,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h5,
3'h5,
3'h3,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h7,
3'h0,
3'h0,
3'h7,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h7,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h7,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h5,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h7,
3'h7,
3'h7,
3'h7,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h7,
3'h7,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h7,
3'h7,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h7,
3'h7,
3'h7,
3'h0,
3'h0,
3'h0,
3'h7,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h5,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h3,
3'h3,
3'h2,
3'h3,
3'h2,
3'h7,
3'h5,
3'h7,
3'h3,
3'h3,
3'h2,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h3,
3'h3,
3'h3,
3'h2,
3'h2,
3'h2,
3'h3,
3'h3,
3'h2,
3'h2,
3'h3,
3'h2,
3'h7,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h7,
3'h7,
3'h3,
3'h3,
3'h3,
3'h2,
3'h7,
3'h7,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h7,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h7,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h2,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h2,
3'h2,
3'h2,
3'h2,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h2,
3'h5,
3'h5,
3'h7,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h7,
3'h7,
3'h7,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h3,
3'h3,
3'h3,
3'h3,
3'h2,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h7,
3'h5,
3'h7,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h7,
3'h7,
3'h3,
3'h3,
3'h3,
3'h7,
3'h7,
3'h7,
3'h7,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h7,
3'h7,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h7,
3'h7,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h7,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h3,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h7,
3'h7,
3'h7,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h3,
3'h3,
3'h2,
3'h2,
3'h2,
3'h3,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h3,
3'h7,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h7,
3'h0,
3'h0,
3'h7,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h7,
3'h5,
3'h5,
3'h3,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h3,
3'h7,
3'h5,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h7,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h2,
3'h2,
3'h2,
3'h2,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h7,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h7,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h3,
3'h3,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h2,
3'h3,
3'h7,
3'h7,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h7,
3'h3,
3'h3,
3'h3,
3'h3,
3'h7,
3'h7,
3'h7,
3'h7,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h7,
3'h7,
3'h7,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h7,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h7,
3'h7,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h7,
3'h7,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h3,
3'h3,
3'h3,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h7,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h7,
3'h3,
3'h3,
3'h3,
3'h7,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h7,
3'h3,
3'h3,
3'h3,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h3,
3'h7,
3'h7,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h7,
3'h7,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h3,
3'h7,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h7,
3'h7,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h3,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h7,
3'h7,
3'h7,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h7,
3'h7,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h7,
3'h3,
3'h7,
3'h7,
3'h7,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h7,
3'h7,
3'h7,
3'h7,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h7,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h2,
3'h2,
3'h3,
3'h2,
3'h2,
3'h2,
3'h2,
3'h3,
3'h2,
3'h2,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h2,
3'h2,
3'h2,
3'h3,
3'h3,
3'h3,
3'h3,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h7,
3'h7,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h7,
3'h7,
3'h3,
3'h3,
3'h3,
3'h3,
3'h5,
3'h5,
3'h7,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h7,
3'h7,
3'h5,
3'h3,
3'h3,
3'h3,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h7,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h7,
3'h7,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h7,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h5,
3'h7,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h7,
3'h7,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h7,
3'h7,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h7,
3'h7,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h7,
3'h7,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h7,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h2,
3'h3,
3'h3,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h7,
3'h7,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h7,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h7,
3'h7,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h7,
3'h3,
3'h2,
3'h3,
3'h3,
3'h3,
3'h3,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h7,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h7,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h7,
3'h7,
3'h7,
3'h7,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h5,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h2,
3'h3,
3'h2,
3'h2,
3'h3,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h2,
3'h3,
3'h3,
3'h3,
3'h7,
3'h7,
3'h7,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h7,
3'h7,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h7,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h7,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h2,
3'h3,
3'h2,
3'h2,
3'h2,
3'h2,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h7,
3'h5,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h7,
3'h7,
3'h7,
3'h7,
3'h2,
3'h3,
3'h3,
3'h2,
3'h2,
3'h3,
3'h3,
3'h3,
3'h7,
3'h7,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h7,
3'h7,
3'h7,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h7,
3'h5,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h7,
3'h7,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h3,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h3,
3'h7,
3'h5,
3'h5,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h5,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h7,
3'h7,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h7,
3'h7,
3'h7,
3'h7,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h7,
3'h7,
3'h7,
3'h0,
3'h0,
3'h0,
3'h0,
3'h7,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h7,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h2,
3'h2,
3'h3,
3'h2,
3'h2,
3'h3,
3'h2,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h3,
3'h5,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h7,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h7,
3'h7,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h7,
3'h7,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h2,
3'h3,
3'h3,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h7,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h7,
3'h7,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h3,
3'h3,
3'h3,
3'h7,
3'h7,
3'h7,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h7,
3'h7,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h3,
3'h2,
3'h3,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h2,
3'h3,
3'h2,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h7,
3'h7,
3'h7,
3'h5,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h7,
3'h7,
3'h3,
3'h3,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h0,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h7,
3'h7,
3'h7,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h5,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h2,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h2,
3'h2,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h2,
3'h3,
3'h5,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h5,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h7,
3'h7,
3'h7,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h5,
3'h7,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h7,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h7,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h2,
3'h3,
3'h3,
3'h3,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h2,
3'h2,
3'h2,
3'h3,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h3,
3'h2,
3'h2,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h7,
3'h5,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h7,
3'h7,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h2,
3'h2,
3'h2,
3'h2,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h5,
3'h7,
3'h7,
3'h7,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h7,
3'h7,
3'h7,
3'h7,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h7,
3'h7,
3'h3,
3'h7,
3'h7,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h7,
3'h7,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h5,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h2,
3'h3,
3'h3,
3'h2,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h5,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h7,
3'h5,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h7,
3'h7,
3'h3,
3'h7,
3'h7,
3'h3,
3'h7,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h7,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h3,
3'h2,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h7,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h2,
3'h2,
3'h2,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h2,
3'h2,
3'h3,
3'h3,
3'h2,
3'h2,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h7,
3'h7,
3'h7,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h7,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h2,
3'h2,
3'h2,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h2,
3'h3,
3'h3,
3'h3,
3'h5,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h0,
3'h0,
3'h7,
3'h7,
3'h7,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h7,
3'h7,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h2,
3'h2,
3'h2,
3'h2,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h7,
3'h7,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h5,
3'h5,
3'h7,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h7,
3'h5,
3'h7,
3'h7,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h7,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h3,
3'h5,
3'h5,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h7,
3'h7,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h2,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h3,
3'h3,
3'h3,
3'h2,
3'h3,
3'h3,
3'h2,
3'h7,
3'h7,
3'h7,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h7,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h2,
3'h2,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h2,
3'h3,
3'h2,
3'h2,
3'h3,
3'h7,
3'h7,
3'h5,
3'h7,
3'h7,
3'h0,
3'h0,
3'h0,
3'h0,
3'h7,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h7,
3'h7,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h2,
3'h3,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h7,
3'h7,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h7,
3'h7,
3'h7,
3'h3,
3'h3,
3'h3,
3'h7,
3'h7,
3'h7,
3'h7,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h7,
3'h7,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h2,
3'h2,
3'h2,
3'h2,
3'h3,
3'h7,
3'h5,
3'h7,
3'h7,
3'h7,
3'h0,
3'h0,
3'h0,
3'h0,
3'h7,
3'h0,
3'h0,
3'h7,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h5,
3'h7,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h2,
3'h2,
3'h3,
3'h3,
3'h3,
3'h5,
3'h2,
3'h3,
3'h3,
3'h3,
3'h5,
3'h5,
3'h7,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h7,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h7,
3'h5,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h7,
3'h3,
3'h2,
3'h2,
3'h2,
3'h3,
3'h7,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h7,
3'h7,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h2,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h5,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h7,
3'h7,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h2,
3'h2,
3'h2,
3'h2,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h7,
3'h7,
3'h7,
3'h0,
3'h0,
3'h7,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h7,
3'h7,
3'h5,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h2,
3'h2,
3'h3,
3'h3,
3'h3,
3'h3,
3'h2,
3'h3,
3'h3,
3'h2,
3'h3,
3'h7,
3'h0,
3'h7,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h7,
3'h7,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h7,
3'h5,
3'h0,
3'h7,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h7,
3'h7,
3'h3,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h7,
3'h7,
3'h7,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h5,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h2,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h2,
3'h3,
3'h3,
3'h2,
3'h3,
3'h3,
3'h7,
3'h5,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h7,
3'h0,
3'h7,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h2,
3'h2,
3'h2,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h2,
3'h2,
3'h3,
3'h2,
3'h3,
3'h3,
3'h3,
3'h2,
3'h3,
3'h3,
3'h3,
3'h7,
3'h7,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h7,
3'h5,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h2,
3'h2,
3'h2,
3'h3,
3'h5,
3'h7,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h7,
3'h7,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h7,
3'h7,
3'h7,
3'h7,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h7,
3'h7,
3'h7,
3'h7,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h5,
3'h7,
3'h3,
3'h3,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h3,
3'h7,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h7,
3'h0,
3'h0,
3'h0,
3'h7,
3'h7,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h5,
3'h7,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h2,
3'h3,
3'h3,
3'h2,
3'h3,
3'h3,
3'h3,
3'h5,
3'h7,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h7,
3'h5,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h2,
3'h2,
3'h2,
3'h2,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h3,
3'h5,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h7,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h7,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h7,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h7,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h7,
3'h7,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h7,
3'h5,
3'h7,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h7,
3'h7,
3'h3,
3'h2,
3'h2,
3'h3,
3'h2,
3'h5,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h7,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h7,
3'h7,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h7,
3'h7,
3'h7,
3'h7,
3'h3,
3'h7,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h7,
3'h3,
3'h3,
3'h7,
3'h7,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h7,
3'h7,
3'h7,
3'h7,
3'h3,
3'h3,
3'h3,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h7,
3'h5,
3'h0,
3'h0,
3'h0,
3'h7,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h7,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h7,
3'h7,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h3,
3'h2,
3'h2,
3'h2,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h2,
3'h3,
3'h3,
3'h3,
3'h7,
3'h7,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h7,
3'h7,
3'h7,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h7,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h7,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h7,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h7,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h7,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h7,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h7,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h7,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h7,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h7,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h7,
3'h7,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h3,
3'h3,
3'h5,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h7,
3'h7,
3'h7,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h7,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h7,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h7,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h7,
3'h5,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h7,
3'h3,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h7,
3'h5,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h7,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h7,
3'h7,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h7,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h7,
3'h0,
3'h0,
3'h0,
3'h7,
3'h5,
3'h7,
3'h3,
3'h3,
3'h3,
3'h2,
3'h3,
3'h3,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h3,
3'h5,
3'h0,
3'h0,
3'h0,
3'h7,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h7,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h7,
3'h7,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h5,
3'h5,
3'h7,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h0,
3'h0,
3'h7,
3'h0,
3'h0,
3'h0,
3'h0,
3'h7,
3'h7,
3'h7,
3'h7,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h7,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h5,
3'h5,
3'h7,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h7,
3'h7,
3'h7,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h7,
3'h5,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h7,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h7,
3'h3,
3'h3,
3'h2,
3'h2,
3'h2,
3'h2,
3'h7,
3'h7,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h7,
3'h7,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h7,
3'h7,
3'h0,
3'h0,
3'h7,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h2,
3'h3,
3'h3,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h3,
3'h7,
3'h7,
3'h0,
3'h0,
3'h0,
3'h0,
3'h7,
3'h7,
3'h7,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h7,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h7,
3'h7,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h7,
3'h7,
3'h0,
3'h0,
3'h0,
3'h0,
3'h7,
3'h7,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h7,
3'h2,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h3,
3'h2,
3'h3,
3'h7,
3'h7,
3'h7,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h7,
3'h7,
3'h7,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h7,
3'h0,
3'h0,
3'h0,
3'h0,
3'h7,
3'h0,
3'h0,
3'h7,
3'h0,
3'h0,
3'h0,
3'h0,
3'h7,
3'h0,
3'h0,
3'h7,
3'h0,
3'h0,
3'h0,
3'h0,
3'h7,
3'h0,
3'h0,
3'h7,
3'h0,
3'h0,
3'h0,
3'h0,
3'h7,
3'h0,
3'h0,
3'h7,
3'h0,
3'h0,
3'h0,
3'h0,
3'h7,
3'h0,
3'h0,
3'h7,
3'h0,
3'h0,
3'h0,
3'h0,
3'h7,
3'h0,
3'h0,
3'h7,
3'h0,
3'h0,
3'h0,
3'h0,
3'h7,
3'h0,
3'h0,
3'h7,
3'h0,
3'h0,
3'h0,
3'h0,
3'h7,
3'h0,
3'h0,
3'h7,
3'h0,
3'h7,
3'h0,
3'h0,
3'h7,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h5,
3'h5,
3'h7,
3'h7,
3'h5,
3'h0,
3'h7,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h7,
3'h0,
3'h0,
3'h7,
3'h0,
3'h0,
3'h7,
3'h0,
3'h7,
3'h0,
3'h0,
3'h7,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h7,
3'h7,
3'h3,
3'h7,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h2,
3'h2,
3'h2,
3'h3,
3'h7,
3'h7,
3'h0,
3'h0,
3'h0,
3'h0,
3'h7,
3'h0,
3'h0,
3'h7,
3'h0,
3'h7,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h7,
3'h0,
3'h0,
3'h0,
3'h0,
3'h7,
3'h0,
3'h7,
3'h7,
3'h7,
3'h7,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h7,
3'h2,
3'h3,
3'h3,
3'h3,
3'h3,
3'h5,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h2,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h3,
3'h7,
3'h7,
3'h7,
3'h0,
3'h0,
3'h7,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h7,
3'h3,
3'h3,
3'h2,
3'h2,
3'h3,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h3,
3'h2,
3'h5,
3'h7,
3'h7,
3'h0,
3'h0,
3'h0,
3'h7,
3'h0,
3'h7,
3'h7,
3'h0,
3'h7,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h7,
3'h7,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h7,
3'h0,
3'h0,
3'h0,
3'h7,
3'h7,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h3,
3'h2,
3'h2,
3'h3,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h7,
3'h5,
3'h7,
3'h5,
3'h0,
3'h7,
3'h0,
3'h0,
3'h0,
3'h0,
3'h7,
3'h0,
3'h7,
3'h0,
3'h0,
3'h7,
3'h0,
3'h7,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h7,
3'h0,
3'h0,
3'h0,
3'h0,
3'h7,
3'h0,
3'h0,
3'h7,
3'h0,
3'h0,
3'h0,
3'h0,
3'h7,
3'h0,
3'h0,
3'h7,
3'h0,
3'h0,
3'h0,
3'h0,
3'h7,
3'h0,
3'h0,
3'h7,
3'h0,
3'h0,
3'h0,
3'h0,
3'h7,
3'h0,
3'h0,
3'h7,
3'h0,
3'h0,
3'h0,
3'h0,
3'h7,
3'h0,
3'h0,
3'h7,
3'h0,
3'h0,
3'h0,
3'h0,
3'h7,
3'h0,
3'h0,
3'h7,
3'h0,
3'h0,
3'h0,
3'h0,
3'h7,
3'h0,
3'h0,
3'h7,
3'h0,
3'h0,
3'h0,
3'h0,
3'h7,
3'h0,
3'h0,
3'h7,
3'h0,
3'h0,
3'h0,
3'h0,
3'h7,
3'h0,
3'h0,
3'h7,
3'h0,
3'h0,
3'h0,
3'h0,
3'h7,
3'h0,
3'h0,
3'h7,
3'h0,
3'h0,
3'h0,
3'h0,
3'h7,
3'h0,
3'h0,
3'h7,
3'h0,
3'h0,
3'h0,
3'h0,
3'h7,
3'h0,
3'h0,
3'h7,
3'h0,
3'h0,
3'h0,
3'h0,
3'h7,
3'h0,
3'h0,
3'h7,
3'h0,
3'h0,
3'h0,
3'h0,
3'h7,
3'h0,
3'h0,
3'h7,
3'h0,
3'h0,
3'h0,
3'h0,
3'h7,
3'h0,
3'h0,
3'h7,
3'h0,
3'h0,
3'h0,
3'h0,
3'h7,
3'h0,
3'h0,
3'h7,
3'h0,
3'h0,
3'h0,
3'h0,
3'h7,
3'h0,
3'h0,
3'h7,
3'h0,
3'h0,
3'h0,
3'h0,
3'h7,
3'h0,
3'h0,
3'h7,
3'h0,
3'h0,
3'h0,
3'h0,
3'h7,
3'h0,
3'h0,
3'h7,
3'h0,
3'h0,
3'h0,
3'h0,
3'h7,
3'h0,
3'h0,
3'h7,
3'h0,
3'h0,
3'h0,
3'h0,
3'h7,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h7,
3'h3,
3'h3,
3'h2,
3'h2,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h3,
3'h2,
3'h2,
3'h3,
3'h2,
3'h2,
3'h3,
3'h3,
3'h3,
3'h5,
3'h7,
3'h7,
3'h0,
3'h0,
3'h7,
3'h0,
3'h0,
3'h7,
3'h0,
3'h7,
3'h0,
3'h0,
3'h0,
3'h0,
3'h7,
3'h0,
3'h0,
3'h7,
3'h0,
3'h0,
3'h0,
3'h0,
3'h7,
3'h0,
3'h0,
3'h7,
3'h0,
3'h0,
3'h0,
3'h0,
3'h7,
3'h0,
3'h0,
3'h7,
3'h0,
3'h0,
3'h0,
3'h0,
3'h7,
3'h0,
3'h0,
3'h0,
3'h7,
3'h0,
3'h0,
3'h7,
3'h0,
3'h7,
3'h0,
3'h0,
3'h7,
3'h0,
3'h0,
3'h7,
3'h0,
3'h7,
3'h0,
3'h0,
3'h7,
3'h0,
3'h0,
3'h7,
3'h0,
3'h7,
3'h0,
3'h0,
3'h7,
3'h0,
3'h0,
3'h7,
3'h0,
3'h7,
3'h0,
3'h0,
3'h7,
3'h0,
3'h0,
3'h7,
3'h0,
3'h7,
3'h0,
3'h0,
3'h7,
3'h0,
3'h0,
3'h7,
3'h0,
3'h7,
3'h0,
3'h0,
3'h7,
3'h0,
3'h0,
3'h7,
3'h0,
3'h7,
3'h0,
3'h0,
3'h7,
3'h0,
3'h0,
3'h7,
3'h0,
3'h7,
3'h7,
3'h0,
3'h7,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h7,
3'h7,
3'h0,
3'h0,
3'h5,
3'h7,
3'h2,
3'h2,
3'h2,
3'h2,
3'h3,
3'h5,
3'h5,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h7,
3'h0,
3'h0,
3'h0,
3'h7,
3'h0,
3'h0,
3'h7,
3'h0,
3'h7,
3'h0,
3'h0,
3'h7,
3'h0,
3'h0,
3'h7,
3'h0,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h7,
3'h7,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h2,
3'h2,
3'h3,
3'h7,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h7,
3'h0,
3'h7,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h7,
3'h0,
3'h7,
3'h0,
3'h7,
3'h7,
3'h7,
3'h7,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h7,
3'h3,
3'h7,
3'h3,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h7,
3'h7,
3'h5,
3'h5,
3'h7,
3'h7,
3'h0,
3'h5,
3'h7,
3'h7,
3'h7,
3'h5,
3'h0,
3'h0,
3'h0,
3'h7,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h7,
3'h3,
3'h3,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h3,
3'h3,
3'h5,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h7,
3'h0,
3'h7,
3'h7,
3'h0,
3'h0,
3'h0,
3'h0,
3'h7,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h7,
3'h0,
3'h0,
3'h0,
3'h7,
3'h7,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h7,
3'h5,
3'h0,
3'h0,
3'h0,
3'h7,
3'h7,
3'h0,
3'h0,
3'h0,
3'h7,
3'h0,
3'h0,
3'h7,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h7,
3'h0,
3'h0,
3'h7,
3'h0,
3'h7,
3'h0,
3'h0,
3'h7,
3'h0,
3'h0,
3'h7,
3'h0,
3'h7,
3'h0,
3'h0,
3'h7,
3'h0,
3'h0,
3'h7,
3'h0,
3'h7,
3'h0,
3'h0,
3'h7,
3'h0,
3'h0,
3'h7,
3'h0,
3'h7,
3'h0,
3'h0,
3'h7,
3'h0,
3'h0,
3'h7,
3'h0,
3'h7,
3'h0,
3'h0,
3'h7,
3'h0,
3'h0,
3'h7,
3'h0,
3'h7,
3'h0,
3'h0,
3'h7,
3'h0,
3'h0,
3'h7,
3'h0,
3'h7,
3'h0,
3'h0,
3'h7,
3'h0,
3'h0,
3'h7,
3'h0,
3'h7,
3'h0,
3'h0,
3'h7,
3'h0,
3'h0,
3'h7,
3'h0,
3'h7,
3'h0,
3'h0,
3'h7,
3'h0,
3'h0,
3'h7,
3'h0,
3'h7,
3'h0,
3'h0,
3'h7,
3'h0,
3'h0,
3'h7,
3'h0,
3'h7,
3'h0,
3'h0,
3'h7,
3'h0,
3'h0,
3'h7,
3'h0,
3'h7,
3'h0,
3'h0,
3'h7,
3'h0,
3'h0,
3'h7,
3'h0,
3'h7,
3'h0,
3'h0,
3'h7,
3'h0,
3'h0,
3'h7,
3'h0,
3'h7,
3'h0,
3'h0,
3'h7,
3'h0,
3'h0,
3'h7,
3'h0,
3'h7,
3'h0,
3'h0,
3'h7,
3'h0,
3'h0,
3'h7,
3'h0,
3'h7,
3'h0,
3'h0,
3'h7,
3'h0,
3'h0,
3'h7,
3'h0,
3'h7,
3'h0,
3'h0,
3'h7,
3'h0,
3'h0,
3'h7,
3'h0,
3'h7,
3'h0,
3'h0,
3'h7,
3'h0,
3'h0,
3'h7,
3'h0,
3'h7,
3'h0,
3'h0,
3'h7,
3'h0,
3'h0,
3'h7,
3'h0,
3'h7,
3'h0,
3'h0,
3'h7,
3'h0,
3'h0,
3'h7,
3'h0,
3'h7,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h7,
3'h7,
3'h0,
3'h5,
3'h5,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h3,
3'h2,
3'h2,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h7,
3'h7,
3'h0,
3'h7,
3'h7,
3'h0,
3'h0,
3'h0,
3'h0,
3'h7,
3'h0,
3'h0,
3'h7,
3'h0,
3'h7,
3'h0,
3'h0,
3'h7,
3'h0,
3'h0,
3'h7,
3'h0,
3'h7,
3'h0,
3'h0,
3'h7,
3'h0,
3'h0,
3'h7,
3'h0,
3'h7,
3'h0,
3'h0,
3'h7,
3'h0,
3'h0,
3'h7,
3'h0,
3'h0,
3'h0,
3'h0,
3'h7,
3'h0,
3'h0,
3'h7,
3'h0,
3'h7,
3'h0,
3'h0,
3'h7,
3'h0,
3'h0,
3'h7,
3'h0,
3'h7,
3'h0,
3'h0,
3'h7,
3'h0,
3'h0,
3'h7,
3'h0,
3'h7,
3'h0,
3'h0,
3'h7,
3'h0,
3'h0,
3'h7,
3'h0,
3'h7,
3'h0,
3'h0,
3'h7,
3'h0,
3'h0,
3'h7,
3'h0,
3'h7,
3'h0,
3'h0,
3'h7,
3'h0,
3'h0,
3'h7,
3'h0,
3'h7,
3'h0,
3'h0,
3'h7,
3'h0,
3'h0,
3'h7,
3'h0,
3'h7,
3'h0,
3'h0,
3'h7,
3'h0,
3'h0,
3'h7,
3'h0,
3'h7,
3'h7,
3'h7,
3'h7,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h7,
3'h7,
3'h7,
3'h3,
3'h3,
3'h3,
3'h2,
3'h2,
3'h2,
3'h2,
3'h3,
3'h3,
3'h7,
3'h7,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h7,
3'h0,
3'h0,
3'h7,
3'h0,
3'h7,
3'h0,
3'h0,
3'h7,
3'h0,
3'h0,
3'h7,
3'h0,
3'h7,
3'h7,
3'h7,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h7,
3'h7,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h2,
3'h2,
3'h2,
3'h2,
3'h3,
3'h5,
3'h7,
3'h0,
3'h0,
3'h7,
3'h0,
3'h7,
3'h7,
3'h0,
3'h0,
3'h0,
3'h0,
3'h7,
3'h0,
3'h7,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h7,
3'h0,
3'h0,
3'h0,
3'h0,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h3,
3'h3,
3'h7,
3'h7,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h5,
3'h7,
3'h7,
3'h7,
3'h5,
3'h7,
3'h5,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h7,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h3,
3'h5,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h0,
3'h0,
3'h7,
3'h7,
3'h7,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h7,
3'h0,
3'h0,
3'h5,
3'h7,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h2,
3'h2,
3'h2,
3'h3,
3'h3,
3'h2,
3'h2,
3'h2,
3'h2,
3'h3,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h7,
3'h7,
3'h7,
3'h7,
3'h0,
3'h7,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h7,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h7,
3'h0,
3'h0,
3'h7,
3'h0,
3'h7,
3'h0,
3'h0,
3'h7,
3'h0,
3'h0,
3'h7,
3'h0,
3'h7,
3'h0,
3'h0,
3'h7,
3'h0,
3'h0,
3'h7,
3'h0,
3'h7,
3'h0,
3'h0,
3'h7,
3'h0,
3'h0,
3'h7,
3'h0,
3'h7,
3'h0,
3'h0,
3'h7,
3'h0,
3'h0,
3'h7,
3'h0,
3'h7,
3'h0,
3'h0,
3'h7,
3'h0,
3'h0,
3'h7,
3'h0,
3'h7,
3'h0,
3'h0,
3'h7,
3'h0,
3'h0,
3'h7,
3'h0,
3'h7,
3'h0,
3'h0,
3'h7,
3'h0,
3'h0,
3'h7,
3'h0,
3'h7,
3'h0,
3'h0,
3'h7,
3'h0,
3'h0,
3'h7,
3'h0,
3'h7,
3'h0,
3'h0,
3'h7,
3'h0,
3'h0,
3'h7,
3'h0,
3'h7,
3'h0,
3'h0,
3'h7,
3'h0,
3'h0,
3'h7,
3'h0,
3'h7,
3'h0,
3'h0,
3'h7,
3'h0,
3'h0,
3'h7,
3'h0,
3'h7,
3'h0,
3'h0,
3'h7,
3'h0,
3'h0,
3'h7,
3'h0,
3'h7,
3'h0,
3'h0,
3'h7,
3'h0,
3'h0,
3'h7,
3'h0,
3'h7,
3'h0,
3'h0,
3'h7,
3'h0,
3'h0,
3'h7,
3'h0,
3'h7,
3'h0,
3'h0,
3'h7,
3'h0,
3'h0,
3'h7,
3'h0,
3'h7,
3'h0,
3'h0,
3'h7,
3'h0,
3'h0,
3'h7,
3'h0,
3'h7,
3'h0,
3'h0,
3'h7,
3'h0,
3'h0,
3'h7,
3'h0,
3'h7,
3'h0,
3'h0,
3'h7,
3'h0,
3'h0,
3'h7,
3'h0,
3'h7,
3'h0,
3'h0,
3'h7,
3'h0,
3'h0,
3'h7,
3'h0,
3'h7,
3'h0,
3'h0,
3'h7,
3'h0,
3'h0,
3'h7,
3'h0,
3'h7,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h7,
3'h5,
3'h2,
3'h3,
3'h3,
3'h2,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h3,
3'h3,
3'h3,
3'h3,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h3,
3'h2,
3'h2,
3'h2,
3'h2,
3'h3,
3'h2,
3'h2,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h7,
3'h7,
3'h7,
3'h7,
3'h0,
3'h0,
3'h0,
3'h0,
3'h7,
3'h0,
3'h0,
3'h7,
3'h0,
3'h7,
3'h0,
3'h0,
3'h7,
3'h0,
3'h0,
3'h7,
3'h0,
3'h7,
3'h0,
3'h0,
3'h7,
3'h0,
3'h0,
3'h7,
3'h0,
3'h7,
3'h0,
3'h0,
3'h7,
3'h0,
3'h0,
3'h7,
3'h0,
3'h0,
3'h0,
3'h7,
3'h0,
3'h0,
3'h0,
3'h0,
3'h7,
3'h0,
3'h0,
3'h7,
3'h0,
3'h0,
3'h0,
3'h0,
3'h7,
3'h0,
3'h0,
3'h7,
3'h0,
3'h0,
3'h0,
3'h0,
3'h7,
3'h0,
3'h0,
3'h7,
3'h0,
3'h0,
3'h0,
3'h0,
3'h7,
3'h0,
3'h0,
3'h7,
3'h0,
3'h0,
3'h0,
3'h0,
3'h7,
3'h0,
3'h0,
3'h7,
3'h0,
3'h0,
3'h0,
3'h0,
3'h7,
3'h0,
3'h0,
3'h7,
3'h0,
3'h0,
3'h0,
3'h0,
3'h7,
3'h0,
3'h0,
3'h7,
3'h0,
3'h0,
3'h0,
3'h0,
3'h7,
3'h0,
3'h7,
3'h7,
3'h0,
3'h7,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h5,
3'h3,
3'h3,
3'h3,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h3,
3'h7,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h7,
3'h0,
3'h0,
3'h0,
3'h0,
3'h7,
3'h0,
3'h0,
3'h7,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h7,
3'h7,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h7,
3'h7,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h3,
3'h5,
3'h5,
3'h0,
3'h7,
3'h7,
3'h0,
3'h7,
3'h0,
3'h0,
3'h7,
3'h0,
3'h0,
3'h7,
3'h0,
3'h0,
3'h0,
3'h0,
3'h7,
3'h0,
3'h0,
3'h7,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h7,
3'h0,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h5,
3'h5,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h3,
3'h3,
3'h3,
3'h7,
3'h3,
3'h7,
3'h3,
3'h7,
3'h5,
3'h7,
3'h5,
3'h7,
3'h7,
3'h5,
3'h5,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h7,
3'h7,
3'h5,
3'h7,
3'h7,
3'h7,
3'h7,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h5,
3'h5,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h3,
3'h7,
3'h5,
3'h5,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h7,
3'h0,
3'h7,
3'h7,
3'h0,
3'h7,
3'h7,
3'h2,
3'h3,
3'h3,
3'h3,
3'h7,
3'h5,
3'h5,
3'h7,
3'h7,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h7,
3'h0,
3'h7,
3'h7,
3'h7,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h7,
3'h7,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h7,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h7,
3'h0,
3'h0,
3'h0,
3'h0,
3'h7,
3'h0,
3'h0,
3'h7,
3'h0,
3'h0,
3'h0,
3'h0,
3'h7,
3'h0,
3'h0,
3'h7,
3'h0,
3'h0,
3'h0,
3'h0,
3'h7,
3'h0,
3'h0,
3'h7,
3'h0,
3'h0,
3'h0,
3'h0,
3'h7,
3'h0,
3'h0,
3'h7,
3'h0,
3'h0,
3'h0,
3'h0,
3'h7,
3'h0,
3'h0,
3'h7,
3'h0,
3'h0,
3'h0,
3'h0,
3'h7,
3'h0,
3'h0,
3'h7,
3'h0,
3'h0,
3'h0,
3'h0,
3'h7,
3'h0,
3'h0,
3'h7,
3'h0,
3'h0,
3'h0,
3'h0,
3'h7,
3'h0,
3'h0,
3'h7,
3'h0,
3'h0,
3'h0,
3'h0,
3'h7,
3'h0,
3'h0,
3'h7,
3'h0,
3'h0,
3'h0,
3'h0,
3'h7,
3'h0,
3'h0,
3'h7,
3'h0,
3'h0,
3'h0,
3'h0,
3'h7,
3'h0,
3'h0,
3'h7,
3'h0,
3'h0,
3'h0,
3'h0,
3'h7,
3'h0,
3'h0,
3'h7,
3'h0,
3'h0,
3'h0,
3'h0,
3'h7,
3'h0,
3'h0,
3'h7,
3'h0,
3'h0,
3'h0,
3'h0,
3'h7,
3'h0,
3'h0,
3'h7,
3'h0,
3'h0,
3'h0,
3'h0,
3'h7,
3'h0,
3'h0,
3'h7,
3'h0,
3'h0,
3'h0,
3'h0,
3'h7,
3'h0,
3'h0,
3'h7,
3'h0,
3'h0,
3'h0,
3'h0,
3'h7,
3'h0,
3'h0,
3'h7,
3'h0,
3'h0,
3'h0,
3'h0,
3'h7,
3'h0,
3'h0,
3'h7,
3'h0,
3'h0,
3'h0,
3'h0,
3'h7,
3'h0,
3'h0,
3'h7,
3'h0,
3'h0,
3'h0,
3'h0,
3'h7,
3'h0,
3'h0,
3'h7,
3'h0,
3'h0,
3'h0,
3'h0,
3'h7,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h7,
3'h7,
3'h5,
3'h3,
3'h3,
3'h3,
3'h2,
3'h3,
3'h2,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h2,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h7,
3'h7,
3'h0,
3'h0,
3'h0,
3'h0,
3'h7,
3'h0,
3'h0,
3'h0,
3'h0,
3'h7,
3'h0,
3'h0,
3'h7,
3'h0,
3'h0,
3'h0,
3'h0,
3'h7,
3'h0,
3'h0,
3'h7,
3'h0,
3'h0,
3'h0,
3'h0,
3'h7,
3'h0,
3'h0,
3'h7,
3'h0,
3'h0,
3'h0,
3'h0,
3'h7,
3'h0,
3'h0,
3'h7,
3'h0,
3'h0,
3'h0,
3'h0,
3'h7,
3'h0,
3'h0,
3'h7,
3'h0,
3'h0,
3'h0,
3'h0,
3'h7,
3'h0,
3'h0,
3'h7,
3'h0,
3'h0,
3'h0,
3'h0,
3'h7,
3'h0,
3'h0,
3'h7,
3'h0,
3'h0,
3'h0,
3'h0,
3'h7,
3'h0,
3'h0,
3'h7,
3'h0,
3'h0,
3'h0,
3'h0,
3'h7,
3'h0,
3'h0,
3'h7,
3'h0,
3'h0,
3'h0,
3'h0,
3'h7,
3'h0,
3'h0,
3'h7,
3'h0,
3'h0,
3'h0,
3'h0,
3'h7,
3'h0,
3'h0,
3'h7,
3'h0,
3'h0,
3'h0,
3'h0,
3'h7,
3'h0,
3'h7,
3'h7,
3'h0,
3'h7,
3'h0,
3'h0,
3'h7,
3'h0,
3'h7,
3'h7,
3'h7,
3'h7,
3'h3,
3'h3,
3'h3,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h3,
3'h7,
3'h0,
3'h7,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h7,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h7,
3'h0,
3'h0,
3'h0,
3'h0,
3'h7,
3'h0,
3'h0,
3'h7,
3'h7,
3'h7,
3'h3,
3'h3,
3'h3,
3'h3,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h7,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h3,
3'h3,
3'h3,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h0,
3'h0,
3'h7,
3'h0,
3'h0,
3'h0,
3'h0,
3'h7,
3'h0,
3'h0,
3'h7,
3'h0,
3'h0,
3'h7,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h7,
3'h0,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h0,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h0,
3'h7,
3'h7,
3'h5,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h7,
3'h7,
3'h7,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h3,
3'h3,
3'h5,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h7,
3'h7,
3'h3,
3'h3,
3'h3,
3'h2,
3'h2,
3'h2,
3'h3,
3'h3,
3'h7,
3'h5,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h7,
3'h0,
3'h7,
3'h7,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h3,
3'h2,
3'h3,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h7,
3'h7,
3'h7,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h7,
3'h0,
3'h7,
3'h7,
3'h0,
3'h7,
3'h0,
3'h0,
3'h7,
3'h0,
3'h0,
3'h0,
3'h0,
3'h7,
3'h0,
3'h0,
3'h7,
3'h0,
3'h0,
3'h0,
3'h0,
3'h7,
3'h0,
3'h0,
3'h7,
3'h0,
3'h0,
3'h0,
3'h0,
3'h7,
3'h0,
3'h0,
3'h7,
3'h0,
3'h0,
3'h0,
3'h0,
3'h7,
3'h0,
3'h0,
3'h7,
3'h0,
3'h0,
3'h0,
3'h0,
3'h7,
3'h0,
3'h0,
3'h7,
3'h0,
3'h0,
3'h0,
3'h0,
3'h7,
3'h0,
3'h0,
3'h7,
3'h0,
3'h0,
3'h0,
3'h0,
3'h7,
3'h0,
3'h0,
3'h7,
3'h0,
3'h0,
3'h0,
3'h0,
3'h7,
3'h0,
3'h0,
3'h7,
3'h0,
3'h0,
3'h0,
3'h0,
3'h7,
3'h0,
3'h0,
3'h7,
3'h0,
3'h0,
3'h0,
3'h0,
3'h7,
3'h0,
3'h0,
3'h7,
3'h0,
3'h0,
3'h0,
3'h0,
3'h7,
3'h0,
3'h0,
3'h7,
3'h0,
3'h0,
3'h0,
3'h0,
3'h7,
3'h0,
3'h0,
3'h7,
3'h0,
3'h0,
3'h0,
3'h0,
3'h7,
3'h0,
3'h0,
3'h7,
3'h0,
3'h0,
3'h0,
3'h0,
3'h7,
3'h0,
3'h0,
3'h7,
3'h0,
3'h0,
3'h0,
3'h0,
3'h7,
3'h0,
3'h0,
3'h7,
3'h0,
3'h0,
3'h0,
3'h0,
3'h7,
3'h0,
3'h0,
3'h7,
3'h0,
3'h0,
3'h0,
3'h0,
3'h7,
3'h0,
3'h0,
3'h7,
3'h0,
3'h0,
3'h0,
3'h0,
3'h7,
3'h0,
3'h0,
3'h7,
3'h0,
3'h0,
3'h0,
3'h0,
3'h7,
3'h0,
3'h0,
3'h7,
3'h0,
3'h0,
3'h0,
3'h0,
3'h7,
3'h0,
3'h0,
3'h7,
3'h0,
3'h0,
3'h0,
3'h0,
3'h7,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h7,
3'h0,
3'h7,
3'h7,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h2,
3'h2,
3'h2,
3'h2,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h7,
3'h7,
3'h0,
3'h0,
3'h0,
3'h0,
3'h7,
3'h0,
3'h0,
3'h0,
3'h0,
3'h7,
3'h0,
3'h0,
3'h7,
3'h0,
3'h0,
3'h0,
3'h0,
3'h7,
3'h0,
3'h0,
3'h7,
3'h0,
3'h0,
3'h0,
3'h0,
3'h7,
3'h0,
3'h0,
3'h7,
3'h0,
3'h0,
3'h0,
3'h0,
3'h7,
3'h0,
3'h0,
3'h0,
3'h7,
3'h0,
3'h0,
3'h7,
3'h0,
3'h7,
3'h0,
3'h0,
3'h7,
3'h0,
3'h0,
3'h7,
3'h0,
3'h7,
3'h0,
3'h0,
3'h7,
3'h0,
3'h0,
3'h7,
3'h0,
3'h7,
3'h0,
3'h0,
3'h7,
3'h0,
3'h0,
3'h7,
3'h0,
3'h7,
3'h0,
3'h0,
3'h7,
3'h0,
3'h0,
3'h7,
3'h0,
3'h7,
3'h0,
3'h0,
3'h7,
3'h0,
3'h0,
3'h7,
3'h0,
3'h7,
3'h0,
3'h0,
3'h7,
3'h0,
3'h0,
3'h7,
3'h0,
3'h7,
3'h0,
3'h0,
3'h7,
3'h0,
3'h0,
3'h7,
3'h0,
3'h0,
3'h0,
3'h0,
3'h7,
3'h0,
3'h0,
3'h7,
3'h0,
3'h7,
3'h7,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h2,
3'h3,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h5,
3'h5,
3'h7,
3'h0,
3'h0,
3'h0,
3'h0,
3'h7,
3'h0,
3'h0,
3'h7,
3'h0,
3'h0,
3'h7,
3'h0,
3'h0,
3'h0,
3'h0,
3'h7,
3'h0,
3'h0,
3'h7,
3'h0,
3'h7,
3'h7,
3'h0,
3'h0,
3'h7,
3'h7,
3'h3,
3'h3,
3'h7,
3'h5,
3'h5,
3'h5,
3'h5,
3'h0,
3'h7,
3'h7,
3'h7,
3'h5,
3'h7,
3'h7,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h7,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h2,
3'h2,
3'h2,
3'h2,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h7,
3'h5,
3'h5,
3'h7,
3'h0,
3'h0,
3'h0,
3'h0,
3'h7,
3'h0,
3'h7,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h7,
3'h0,
3'h0,
3'h0,
3'h7,
3'h0,
3'h0,
3'h7,
3'h0,
3'h0,
3'h7,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h7,
3'h0,
3'h0,
3'h0,
3'h0,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h0,
3'h7,
3'h7,
3'h0,
3'h7,
3'h7,
3'h7,
3'h7,
3'h0,
3'h7,
3'h7,
3'h0,
3'h7,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h7,
3'h7,
3'h7,
3'h0,
3'h0,
3'h0,
3'h0,
3'h7,
3'h2,
3'h2,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h2,
3'h2,
3'h2,
3'h2,
3'h3,
3'h2,
3'h3,
3'h3,
3'h2,
3'h2,
3'h7,
3'h5,
3'h7,
3'h0,
3'h0,
3'h0,
3'h0,
3'h7,
3'h5,
3'h7,
3'h3,
3'h3,
3'h3,
3'h3,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h7,
3'h0,
3'h7,
3'h0,
3'h7,
3'h0,
3'h7,
3'h0,
3'h0,
3'h7,
3'h5,
3'h7,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h3,
3'h3,
3'h3,
3'h3,
3'h2,
3'h2,
3'h2,
3'h2,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h2,
3'h3,
3'h3,
3'h3,
3'h3,
3'h7,
3'h7,
3'h5,
3'h3,
3'h0,
3'h0,
3'h7,
3'h0,
3'h0,
3'h0,
3'h0,
3'h7,
3'h0,
3'h0,
3'h7,
3'h0,
3'h0,
3'h0,
3'h0,
3'h7,
3'h0,
3'h0,
3'h7,
3'h0,
3'h7,
3'h0,
3'h0,
3'h7,
3'h0,
3'h0,
3'h7,
3'h0,
3'h7,
3'h0,
3'h0,
3'h7,
3'h0,
3'h0,
3'h7,
3'h0,
3'h7,
3'h0,
3'h0,
3'h7,
3'h0,
3'h0,
3'h7,
3'h0,
3'h7,
3'h0,
3'h0,
3'h7,
3'h0,
3'h0,
3'h7,
3'h0,
3'h7,
3'h0,
3'h0,
3'h7,
3'h0,
3'h0,
3'h7,
3'h0,
3'h7,
3'h0,
3'h0,
3'h7,
3'h0,
3'h0,
3'h7,
3'h0,
3'h7,
3'h0,
3'h0,
3'h7,
3'h0,
3'h0,
3'h7,
3'h0,
3'h7,
3'h0,
3'h0,
3'h7,
3'h0,
3'h0,
3'h7,
3'h0,
3'h7,
3'h0,
3'h0,
3'h7,
3'h0,
3'h0,
3'h7,
3'h0,
3'h7,
3'h0,
3'h0,
3'h7,
3'h0,
3'h0,
3'h7,
3'h0,
3'h7,
3'h0,
3'h0,
3'h7,
3'h0,
3'h0,
3'h7,
3'h0,
3'h7,
3'h0,
3'h0,
3'h7,
3'h0,
3'h0,
3'h7,
3'h0,
3'h7,
3'h0,
3'h0,
3'h7,
3'h0,
3'h0,
3'h7,
3'h0,
3'h7,
3'h0,
3'h0,
3'h7,
3'h0,
3'h0,
3'h7,
3'h0,
3'h7,
3'h0,
3'h0,
3'h7,
3'h0,
3'h0,
3'h7,
3'h0,
3'h7,
3'h0,
3'h0,
3'h7,
3'h0,
3'h0,
3'h7,
3'h0,
3'h7,
3'h0,
3'h0,
3'h7,
3'h0,
3'h0,
3'h7,
3'h0,
3'h7,
3'h0,
3'h0,
3'h7,
3'h0,
3'h0,
3'h7,
3'h0,
3'h7,
3'h0,
3'h0,
3'h7,
3'h0,
3'h0,
3'h7,
3'h0,
3'h7,
3'h0,
3'h0,
3'h7,
3'h0,
3'h0,
3'h7,
3'h0,
3'h7,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h7,
3'h0,
3'h7,
3'h3,
3'h3,
3'h2,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h2,
3'h2,
3'h2,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h7,
3'h7,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h7,
3'h0,
3'h0,
3'h7,
3'h0,
3'h7,
3'h0,
3'h0,
3'h7,
3'h0,
3'h0,
3'h7,
3'h0,
3'h7,
3'h0,
3'h0,
3'h7,
3'h0,
3'h0,
3'h7,
3'h0,
3'h7,
3'h0,
3'h0,
3'h7,
3'h0,
3'h0,
3'h7,
3'h0,
3'h0,
3'h0,
3'h0,
3'h7,
3'h0,
3'h0,
3'h7,
3'h0,
3'h0,
3'h0,
3'h0,
3'h7,
3'h0,
3'h0,
3'h7,
3'h0,
3'h0,
3'h0,
3'h0,
3'h7,
3'h0,
3'h0,
3'h7,
3'h0,
3'h0,
3'h0,
3'h0,
3'h7,
3'h0,
3'h0,
3'h7,
3'h0,
3'h0,
3'h0,
3'h0,
3'h7,
3'h0,
3'h0,
3'h7,
3'h0,
3'h0,
3'h0,
3'h0,
3'h7,
3'h0,
3'h0,
3'h7,
3'h0,
3'h0,
3'h0,
3'h0,
3'h7,
3'h0,
3'h0,
3'h7,
3'h0,
3'h0,
3'h0,
3'h0,
3'h7,
3'h0,
3'h0,
3'h7,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h7,
3'h7,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h3,
3'h3,
3'h7,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h7,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h7,
3'h0,
3'h0,
3'h7,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h7,
3'h7,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h2,
3'h3,
3'h2,
3'h2,
3'h5,
3'h2,
3'h7,
3'h0,
3'h0,
3'h0,
3'h0,
3'h7,
3'h7,
3'h0,
3'h0,
3'h0,
3'h7,
3'h0,
3'h0,
3'h7,
3'h0,
3'h0,
3'h0,
3'h7,
3'h7,
3'h7,
3'h7,
3'h0,
3'h0,
3'h0,
3'h7,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h7,
3'h7,
3'h7,
3'h7,
3'h0,
3'h7,
3'h0,
3'h7,
3'h7,
3'h0,
3'h7,
3'h0,
3'h0,
3'h7,
3'h7,
3'h0,
3'h7,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h7,
3'h7,
3'h7,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h7,
3'h0,
3'h0,
3'h7,
3'h2,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h2,
3'h2,
3'h2,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h2,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h2,
3'h2,
3'h2,
3'h3,
3'h3,
3'h7,
3'h0,
3'h7,
3'h0,
3'h7,
3'h7,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h2,
3'h3,
3'h2,
3'h3,
3'h2,
3'h3,
3'h5,
3'h0,
3'h0,
3'h0,
3'h7,
3'h0,
3'h7,
3'h0,
3'h0,
3'h7,
3'h5,
3'h7,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h2,
3'h2,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h5,
3'h7,
3'h0,
3'h0,
3'h7,
3'h0,
3'h0,
3'h0,
3'h0,
3'h7,
3'h0,
3'h0,
3'h7,
3'h0,
3'h0,
3'h0,
3'h0,
3'h7,
3'h0,
3'h0,
3'h7,
3'h0,
3'h0,
3'h0,
3'h0,
3'h7,
3'h0,
3'h0,
3'h7,
3'h0,
3'h0,
3'h0,
3'h0,
3'h7,
3'h0,
3'h0,
3'h7,
3'h0,
3'h0,
3'h0,
3'h0,
3'h7,
3'h0,
3'h0,
3'h7,
3'h0,
3'h0,
3'h0,
3'h0,
3'h7,
3'h0,
3'h0,
3'h7,
3'h0,
3'h0,
3'h0,
3'h0,
3'h7,
3'h0,
3'h0,
3'h7,
3'h0,
3'h0,
3'h0,
3'h0,
3'h7,
3'h0,
3'h0,
3'h7,
3'h0,
3'h0,
3'h0,
3'h0,
3'h7,
3'h0,
3'h0,
3'h7,
3'h0,
3'h0,
3'h0,
3'h0,
3'h7,
3'h0,
3'h0,
3'h7,
3'h0,
3'h0,
3'h0,
3'h0,
3'h7,
3'h0,
3'h0,
3'h7,
3'h0,
3'h0,
3'h0,
3'h0,
3'h7,
3'h0,
3'h0,
3'h7,
3'h0,
3'h0,
3'h0,
3'h0,
3'h7,
3'h0,
3'h0,
3'h7,
3'h0,
3'h0,
3'h0,
3'h0,
3'h7,
3'h0,
3'h0,
3'h7,
3'h0,
3'h0,
3'h0,
3'h0,
3'h7,
3'h0,
3'h0,
3'h7,
3'h0,
3'h0,
3'h0,
3'h0,
3'h7,
3'h0,
3'h0,
3'h7,
3'h0,
3'h0,
3'h0,
3'h0,
3'h7,
3'h0,
3'h0,
3'h7,
3'h0,
3'h0,
3'h0,
3'h0,
3'h7,
3'h0,
3'h0,
3'h7,
3'h0,
3'h0,
3'h0,
3'h0,
3'h7,
3'h0,
3'h0,
3'h7,
3'h0,
3'h0,
3'h0,
3'h0,
3'h7,
3'h0,
3'h0,
3'h7,
3'h0,
3'h0,
3'h0,
3'h0,
3'h7,
3'h0,
3'h0,
3'h7,
3'h0,
3'h0,
3'h0,
3'h0,
3'h7,
3'h0,
3'h0,
3'h7,
3'h0,
3'h0,
3'h7,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h7,
3'h7,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h2,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h5,
3'h5,
3'h7,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h7,
3'h0,
3'h0,
3'h7,
3'h0,
3'h0,
3'h0,
3'h0,
3'h7,
3'h0,
3'h0,
3'h7,
3'h0,
3'h0,
3'h0,
3'h0,
3'h7,
3'h0,
3'h0,
3'h7,
3'h0,
3'h0,
3'h0,
3'h0,
3'h7,
3'h0,
3'h0,
3'h7,
3'h0,
3'h0,
3'h0,
3'h7,
3'h0,
3'h0,
3'h0,
3'h0,
3'h7,
3'h0,
3'h0,
3'h7,
3'h0,
3'h0,
3'h0,
3'h0,
3'h7,
3'h0,
3'h0,
3'h7,
3'h0,
3'h0,
3'h0,
3'h0,
3'h7,
3'h0,
3'h0,
3'h7,
3'h0,
3'h0,
3'h0,
3'h0,
3'h7,
3'h0,
3'h0,
3'h7,
3'h0,
3'h0,
3'h0,
3'h0,
3'h7,
3'h0,
3'h0,
3'h7,
3'h0,
3'h0,
3'h0,
3'h0,
3'h7,
3'h0,
3'h0,
3'h7,
3'h0,
3'h0,
3'h0,
3'h0,
3'h7,
3'h0,
3'h0,
3'h7,
3'h0,
3'h0,
3'h0,
3'h0,
3'h7,
3'h0,
3'h0,
3'h0,
3'h0,
3'h7,
3'h7,
3'h7,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h7,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h7,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h7,
3'h0,
3'h7,
3'h7,
3'h0,
3'h7,
3'h0,
3'h0,
3'h0,
3'h7,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h7,
3'h7,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h2,
3'h3,
3'h2,
3'h2,
3'h3,
3'h2,
3'h3,
3'h7,
3'h7,
3'h0,
3'h7,
3'h0,
3'h0,
3'h7,
3'h0,
3'h0,
3'h7,
3'h0,
3'h7,
3'h7,
3'h0,
3'h0,
3'h0,
3'h7,
3'h0,
3'h0,
3'h7,
3'h0,
3'h0,
3'h7,
3'h0,
3'h7,
3'h0,
3'h0,
3'h7,
3'h0,
3'h7,
3'h7,
3'h0,
3'h0,
3'h0,
3'h0,
3'h7,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h7,
3'h0,
3'h7,
3'h0,
3'h0,
3'h7,
3'h0,
3'h0,
3'h7,
3'h0,
3'h7,
3'h0,
3'h0,
3'h7,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h7,
3'h0,
3'h0,
3'h0,
3'h0,
3'h7,
3'h0,
3'h7,
3'h0,
3'h0,
3'h0,
3'h0,
3'h7,
3'h7,
3'h0,
3'h7,
3'h7,
3'h7,
3'h7,
3'h3,
3'h3,
3'h3,
3'h2,
3'h3,
3'h3,
3'h3,
3'h3,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h3,
3'h3,
3'h3,
3'h3,
3'h2,
3'h3,
3'h3,
3'h3,
3'h2,
3'h3,
3'h2,
3'h3,
3'h3,
3'h2,
3'h2,
3'h2,
3'h2,
3'h3,
3'h7,
3'h0,
3'h0,
3'h7,
3'h7,
3'h3,
3'h3,
3'h2,
3'h3,
3'h3,
3'h3,
3'h2,
3'h3,
3'h2,
3'h3,
3'h2,
3'h2,
3'h5,
3'h7,
3'h7,
3'h0,
3'h0,
3'h7,
3'h0,
3'h0,
3'h0,
3'h0,
3'h7,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h2,
3'h2,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h2,
3'h2,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h7,
3'h7,
3'h7,
3'h0,
3'h7,
3'h7,
3'h0,
3'h7,
3'h0,
3'h0,
3'h7,
3'h0,
3'h0,
3'h7,
3'h0,
3'h7,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h7,
3'h0,
3'h0,
3'h0,
3'h0,
3'h7,
3'h0,
3'h0,
3'h7,
3'h0,
3'h0,
3'h0,
3'h0,
3'h7,
3'h0,
3'h0,
3'h7,
3'h0,
3'h0,
3'h0,
3'h0,
3'h7,
3'h0,
3'h0,
3'h7,
3'h0,
3'h0,
3'h0,
3'h0,
3'h7,
3'h0,
3'h0,
3'h7,
3'h0,
3'h7,
3'h0,
3'h0,
3'h7,
3'h0,
3'h0,
3'h7,
3'h0,
3'h0,
3'h0,
3'h0,
3'h7,
3'h0,
3'h0,
3'h7,
3'h0,
3'h0,
3'h0,
3'h0,
3'h7,
3'h0,
3'h0,
3'h7,
3'h0,
3'h0,
3'h0,
3'h0,
3'h7,
3'h0,
3'h0,
3'h7,
3'h0,
3'h0,
3'h0,
3'h0,
3'h7,
3'h0,
3'h0,
3'h7,
3'h0,
3'h0,
3'h0,
3'h0,
3'h7,
3'h0,
3'h0,
3'h7,
3'h0,
3'h0,
3'h0,
3'h0,
3'h7,
3'h0,
3'h0,
3'h7,
3'h0,
3'h0,
3'h0,
3'h0,
3'h7,
3'h0,
3'h0,
3'h7,
3'h0,
3'h0,
3'h0,
3'h0,
3'h7,
3'h0,
3'h0,
3'h7,
3'h0,
3'h0,
3'h0,
3'h0,
3'h7,
3'h0,
3'h0,
3'h7,
3'h0,
3'h0,
3'h0,
3'h0,
3'h7,
3'h0,
3'h0,
3'h7,
3'h0,
3'h0,
3'h0,
3'h0,
3'h7,
3'h0,
3'h0,
3'h7,
3'h0,
3'h0,
3'h0,
3'h0,
3'h7,
3'h0,
3'h0,
3'h7,
3'h0,
3'h0,
3'h0,
3'h0,
3'h7,
3'h0,
3'h0,
3'h7,
3'h0,
3'h0,
3'h0,
3'h0,
3'h7,
3'h0,
3'h0,
3'h7,
3'h0,
3'h0,
3'h0,
3'h0,
3'h7,
3'h0,
3'h0,
3'h7,
3'h0,
3'h7,
3'h7,
3'h0,
3'h7,
3'h0,
3'h0,
3'h0,
3'h0,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h0,
3'h0,
3'h0,
3'h7,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h2,
3'h3,
3'h3,
3'h3,
3'h5,
3'h5,
3'h5,
3'h7,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h7,
3'h0,
3'h0,
3'h0,
3'h0,
3'h7,
3'h0,
3'h0,
3'h7,
3'h0,
3'h0,
3'h0,
3'h0,
3'h7,
3'h0,
3'h0,
3'h7,
3'h0,
3'h0,
3'h0,
3'h0,
3'h7,
3'h0,
3'h0,
3'h7,
3'h0,
3'h0,
3'h0,
3'h0,
3'h7,
3'h0,
3'h0,
3'h7,
3'h0,
3'h0,
3'h0,
3'h0,
3'h7,
3'h0,
3'h0,
3'h0,
3'h0,
3'h7,
3'h0,
3'h0,
3'h0,
3'h0,
3'h7,
3'h7,
3'h0,
3'h0,
3'h0,
3'h0,
3'h7,
3'h7,
3'h0,
3'h0,
3'h7,
3'h7,
3'h7,
3'h0,
3'h0,
3'h7,
3'h7,
3'h7,
3'h0,
3'h0,
3'h0,
3'h0,
3'h7,
3'h7,
3'h0,
3'h0,
3'h7,
3'h7,
3'h7,
3'h0,
3'h0,
3'h7,
3'h0,
3'h7,
3'h0,
3'h0,
3'h0,
3'h0,
3'h7,
3'h0,
3'h0,
3'h0,
3'h7,
3'h7,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h7,
3'h7,
3'h7,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h3,
3'h3,
3'h7,
3'h7,
3'h7,
3'h0,
3'h0,
3'h0,
3'h0,
3'h7,
3'h0,
3'h0,
3'h0,
3'h7,
3'h7,
3'h0,
3'h0,
3'h0,
3'h7,
3'h7,
3'h7,
3'h0,
3'h0,
3'h0,
3'h0,
3'h7,
3'h7,
3'h0,
3'h0,
3'h7,
3'h7,
3'h7,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h7,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h7,
3'h5,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h7,
3'h0,
3'h0,
3'h7,
3'h7,
3'h0,
3'h0,
3'h7,
3'h7,
3'h7,
3'h7,
3'h0,
3'h0,
3'h7,
3'h7,
3'h7,
3'h0,
3'h0,
3'h7,
3'h7,
3'h7,
3'h0,
3'h0,
3'h7,
3'h0,
3'h7,
3'h0,
3'h0,
3'h0,
3'h7,
3'h7,
3'h7,
3'h0,
3'h0,
3'h7,
3'h7,
3'h7,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h7,
3'h0,
3'h0,
3'h0,
3'h7,
3'h7,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h7,
3'h0,
3'h0,
3'h0,
3'h0,
3'h7,
3'h0,
3'h0,
3'h0,
3'h7,
3'h7,
3'h0,
3'h7,
3'h3,
3'h3,
3'h3,
3'h2,
3'h3,
3'h3,
3'h3,
3'h3,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h2,
3'h2,
3'h2,
3'h2,
3'h3,
3'h2,
3'h2,
3'h5,
3'h5,
3'h7,
3'h7,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h7,
3'h0,
3'h0,
3'h0,
3'h7,
3'h0,
3'h0,
3'h0,
3'h7,
3'h7,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h7,
3'h5,
3'h0,
3'h0,
3'h7,
3'h7,
3'h7,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h7,
3'h7,
3'h7,
3'h0,
3'h0,
3'h0,
3'h7,
3'h7,
3'h0,
3'h0,
3'h0,
3'h0,
3'h7,
3'h7,
3'h0,
3'h0,
3'h7,
3'h7,
3'h7,
3'h0,
3'h0,
3'h0,
3'h0,
3'h7,
3'h0,
3'h0,
3'h0,
3'h0,
3'h7,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h7,
3'h7,
3'h7,
3'h0,
3'h0,
3'h7,
3'h7,
3'h7,
3'h0,
3'h0,
3'h0,
3'h7,
3'h0,
3'h0,
3'h0,
3'h0,
3'h7,
3'h7,
3'h0,
3'h0,
3'h0,
3'h0,
3'h7,
3'h7,
3'h0,
3'h0,
3'h7,
3'h7,
3'h7,
3'h0,
3'h0,
3'h7,
3'h7,
3'h7,
3'h0,
3'h0,
3'h0,
3'h0,
3'h7,
3'h7,
3'h0,
3'h0,
3'h7,
3'h7,
3'h7,
3'h0,
3'h0,
3'h7,
3'h7,
3'h7,
3'h0,
3'h0,
3'h0,
3'h0,
3'h7,
3'h7,
3'h0,
3'h0,
3'h7,
3'h7,
3'h7,
3'h0,
3'h0,
3'h7,
3'h7,
3'h7,
3'h0,
3'h0,
3'h0,
3'h0,
3'h7,
3'h7,
3'h0,
3'h0,
3'h7,
3'h7,
3'h7,
3'h0,
3'h0,
3'h7,
3'h7,
3'h7,
3'h7,
3'h0,
3'h0,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h0,
3'h0,
3'h0,
3'h0,
3'h7,
3'h7,
3'h0,
3'h0,
3'h0,
3'h7,
3'h7,
3'h0,
3'h0,
3'h7,
3'h7,
3'h7,
3'h7,
3'h0,
3'h0,
3'h7,
3'h7,
3'h7,
3'h0,
3'h0,
3'h0,
3'h7,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h7,
3'h0,
3'h0,
3'h0,
3'h7,
3'h7,
3'h0,
3'h0,
3'h0,
3'h7,
3'h7,
3'h7,
3'h0,
3'h0,
3'h0,
3'h0,
3'h7,
3'h0,
3'h0,
3'h7,
3'h3,
3'h3,
3'h3,
3'h3,
3'h7,
3'h5,
3'h5,
3'h5,
3'h5,
3'h7,
3'h7,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h2,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h7,
3'h5,
3'h5,
3'h5,
3'h7,
3'h7,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h7,
3'h0,
3'h0,
3'h0,
3'h0,
3'h7,
3'h7,
3'h0,
3'h0,
3'h7,
3'h7,
3'h7,
3'h0,
3'h0,
3'h7,
3'h7,
3'h7,
3'h0,
3'h0,
3'h0,
3'h0,
3'h7,
3'h7,
3'h0,
3'h0,
3'h7,
3'h7,
3'h7,
3'h0,
3'h0,
3'h7,
3'h7,
3'h7,
3'h7,
3'h0,
3'h0,
3'h7,
3'h7,
3'h7,
3'h0,
3'h0,
3'h7,
3'h7,
3'h7,
3'h0,
3'h0,
3'h7,
3'h7,
3'h7,
3'h7,
3'h0,
3'h0,
3'h7,
3'h7,
3'h7,
3'h0,
3'h0,
3'h7,
3'h7,
3'h7,
3'h0,
3'h0,
3'h7,
3'h7,
3'h7,
3'h7,
3'h0,
3'h0,
3'h7,
3'h7,
3'h7,
3'h0,
3'h0,
3'h7,
3'h7,
3'h7,
3'h0,
3'h0,
3'h7,
3'h7,
3'h7,
3'h7,
3'h0,
3'h0,
3'h7,
3'h7,
3'h7,
3'h0,
3'h7,
3'h7,
3'h7,
3'h7,
3'h0,
3'h0,
3'h0,
3'h0,
3'h7,
3'h7,
3'h7,
3'h7,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h3,
3'h7,
3'h7,
3'h0,
3'h7,
3'h0,
3'h7,
3'h7,
3'h7,
3'h0,
3'h0,
3'h7,
3'h0,
3'h0,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h0,
3'h0,
3'h0,
3'h7,
3'h7,
3'h7,
3'h0,
3'h0,
3'h7,
3'h7,
3'h7,
3'h0,
3'h7,
3'h7,
3'h7,
3'h0,
3'h0,
3'h0,
3'h0,
3'h7,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h3,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h0,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h0,
3'h0,
3'h7,
3'h7,
3'h7,
3'h0,
3'h0,
3'h7,
3'h7,
3'h7,
3'h0,
3'h0,
3'h7,
3'h7,
3'h7,
3'h7,
3'h0,
3'h0,
3'h7,
3'h7,
3'h7,
3'h0,
3'h0,
3'h7,
3'h7,
3'h7,
3'h0,
3'h0,
3'h7,
3'h7,
3'h7,
3'h0,
3'h0,
3'h0,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h0,
3'h0,
3'h0,
3'h0,
3'h7,
3'h0,
3'h0,
3'h0,
3'h7,
3'h7,
3'h7,
3'h0,
3'h0,
3'h7,
3'h7,
3'h7,
3'h0,
3'h0,
3'h7,
3'h0,
3'h0,
3'h7,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h7,
3'h7,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h2,
3'h2,
3'h2,
3'h2,
3'h3,
3'h3,
3'h3,
3'h7,
3'h7,
3'h7,
3'h7,
3'h0,
3'h0,
3'h7,
3'h5,
3'h5,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h2,
3'h2,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h7,
3'h7,
3'h7,
3'h0,
3'h0,
3'h7,
3'h7,
3'h7,
3'h7,
3'h0,
3'h0,
3'h7,
3'h7,
3'h7,
3'h0,
3'h0,
3'h7,
3'h7,
3'h7,
3'h0,
3'h0,
3'h7,
3'h7,
3'h7,
3'h7,
3'h0,
3'h0,
3'h7,
3'h7,
3'h7,
3'h0,
3'h0,
3'h0,
3'h7,
3'h0,
3'h0,
3'h0,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h0,
3'h0,
3'h0,
3'h7,
3'h7,
3'h0,
3'h0,
3'h7,
3'h7,
3'h7,
3'h7,
3'h0,
3'h0,
3'h7,
3'h7,
3'h7,
3'h0,
3'h0,
3'h7,
3'h7,
3'h7,
3'h0,
3'h0,
3'h7,
3'h7,
3'h7,
3'h7,
3'h0,
3'h0,
3'h7,
3'h7,
3'h7,
3'h0,
3'h0,
3'h7,
3'h7,
3'h7,
3'h0,
3'h0,
3'h7,
3'h7,
3'h7,
3'h7,
3'h0,
3'h0,
3'h7,
3'h7,
3'h7,
3'h0,
3'h0,
3'h7,
3'h7,
3'h7,
3'h0,
3'h0,
3'h7,
3'h7,
3'h7,
3'h7,
3'h0,
3'h0,
3'h7,
3'h7,
3'h7,
3'h0,
3'h0,
3'h7,
3'h7,
3'h7,
3'h0,
3'h0,
3'h7,
3'h7,
3'h7,
3'h7,
3'h0,
3'h0,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h0,
3'h0,
3'h7,
3'h7,
3'h7,
3'h0,
3'h0,
3'h7,
3'h7,
3'h7,
3'h0,
3'h0,
3'h7,
3'h7,
3'h7,
3'h7,
3'h0,
3'h0,
3'h7,
3'h7,
3'h7,
3'h0,
3'h0,
3'h0,
3'h7,
3'h7,
3'h0,
3'h0,
3'h7,
3'h0,
3'h7,
3'h0,
3'h0,
3'h0,
3'h7,
3'h7,
3'h7,
3'h0,
3'h0,
3'h7,
3'h7,
3'h7,
3'h7,
3'h0,
3'h0,
3'h0,
3'h7,
3'h7,
3'h7,
3'h3,
3'h3,
3'h3,
3'h2,
3'h2,
3'h3,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h0,
3'h0,
3'h0,
3'h7,
3'h7,
3'h7,
3'h0,
3'h0,
3'h7,
3'h7,
3'h7,
3'h0,
3'h0,
3'h7,
3'h7,
3'h7,
3'h0,
3'h0,
3'h7,
3'h7,
3'h7,
3'h7,
3'h0,
3'h0,
3'h7,
3'h7,
3'h7,
3'h0,
3'h0,
3'h7,
3'h7,
3'h7,
3'h0,
3'h0,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h0,
3'h7,
3'h7,
3'h7,
3'h7,
3'h0,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h0,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h0,
3'h7,
3'h7,
3'h7,
3'h7,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h7,
3'h5,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h0,
3'h0,
3'h0,
3'h7,
3'h7,
3'h0,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h0,
3'h0,
3'h7,
3'h7,
3'h7,
3'h7,
3'h0,
3'h0,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h0,
3'h7,
3'h7,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h3,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h0,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h0,
3'h7,
3'h7,
3'h7,
3'h7,
3'h0,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h0,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h0,
3'h7,
3'h7,
3'h0,
3'h7,
3'h7,
3'h3,
3'h2,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h2,
3'h2,
3'h2,
3'h3,
3'h2,
3'h2,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h2,
3'h2,
3'h2,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h5,
3'h7,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h0,
3'h0,
3'h0,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h0,
3'h0,
3'h7,
3'h7,
3'h7,
3'h0,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h0,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h0,
3'h7,
3'h7,
3'h7,
3'h7,
3'h0,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h0,
3'h0,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h7,
3'h7,
3'h7,
3'h0,
3'h0,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h0,
3'h0,
3'h7,
3'h3,
3'h3,
3'h3,
3'h3,
3'h2,
3'h2,
3'h2,
3'h2,
3'h3,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h7,
3'h7,
3'h7,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h0,
3'h0,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h2,
3'h3,
3'h3,
3'h3,
3'h3,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h3,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h5,
3'h0,
3'h7,
3'h7,
3'h0,
3'h0,
3'h7,
3'h7,
3'h0,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h0,
3'h7,
3'h7,
3'h0,
3'h0,
3'h7,
3'h7,
3'h0,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h3,
3'h3,
3'h7,
3'h7,
3'h7,
3'h7,
3'h0,
3'h0,
3'h7,
3'h7,
3'h7,
3'h0,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h0,
3'h7,
3'h7,
3'h7,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h2,
3'h3,
3'h3,
3'h3,
3'h3,
3'h2,
3'h2,
3'h2,
3'h7,
3'h7,
3'h5,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h7,
3'h7,
3'h7,
3'h7,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h0,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h0,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h0,
3'h0,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h0,
3'h0,
3'h0,
3'h7,
3'h7,
3'h7,
3'h7,
3'h0,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h0,
3'h7,
3'h0,
3'h0,
3'h0,
3'h7,
3'h7,
3'h7,
3'h7,
3'h0,
3'h0,
3'h7,
3'h7,
3'h0,
3'h0,
3'h7,
3'h7,
3'h7,
3'h3,
3'h3,
3'h3,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h7,
3'h7,
3'h7,
3'h7,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h3,
3'h3,
3'h3,
3'h3,
3'h2,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h2,
3'h3,
3'h3,
3'h3,
3'h3,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h5,
3'h5,
3'h7,
3'h7,
3'h0,
3'h0,
3'h0,
3'h0,
3'h7,
3'h0,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h5,
3'h5,
3'h5,
3'h7,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h7,
3'h7,
3'h0,
3'h7,
3'h7,
3'h0,
3'h0,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h0,
3'h7,
3'h7,
3'h7,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h7,
3'h7,
3'h7,
3'h0,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h0,
3'h0,
3'h7,
3'h0,
3'h7,
3'h7,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h2,
3'h2,
3'h2,
3'h3,
3'h5,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h7,
3'h7,
3'h7,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h7,
3'h7,
3'h7,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h0,
3'h0,
3'h0,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h0,
3'h0,
3'h0,
3'h0,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h0,
3'h0,
3'h0,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h0,
3'h0,
3'h0,
3'h7,
3'h7,
3'h7,
3'h7,
3'h5,
3'h5,
3'h7,
3'h7,
3'h0,
3'h7,
3'h7,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h7,
3'h7,
3'h7,
3'h7,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h0,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h5,
3'h7,
3'h3,
3'h3,
3'h3,
3'h3,
3'h2,
3'h3,
3'h3,
3'h3,
3'h3,
3'h2,
3'h2,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h2,
3'h2,
3'h3,
3'h3,
3'h3,
3'h3,
3'h2,
3'h2,
3'h2,
3'h3,
3'h3,
3'h7,
3'h5,
3'h0,
3'h7,
3'h0,
3'h0,
3'h0,
3'h0,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h0,
3'h7,
3'h7,
3'h7,
3'h7,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h7,
3'h7,
3'h7,
3'h5,
3'h5,
3'h5,
3'h5,
3'h7,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h2,
3'h2,
3'h3,
3'h3,
3'h2,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h7,
3'h7,
3'h7,
3'h7,
3'h0,
3'h0,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h0,
3'h7,
3'h7,
3'h7,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h7,
3'h7,
3'h0,
3'h0,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h0,
3'h7,
3'h7,
3'h0,
3'h0,
3'h0,
3'h0,
3'h7,
3'h7,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h2,
3'h2,
3'h2,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h3,
3'h3,
3'h3,
3'h2,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h2,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h2,
3'h3,
3'h3,
3'h7,
3'h7,
3'h0,
3'h0,
3'h7,
3'h7,
3'h7,
3'h7,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h7,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h7,
3'h7,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h0,
3'h7,
3'h0,
3'h0,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h0,
3'h0,
3'h0,
3'h0,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h0,
3'h0,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h0,
3'h7,
3'h7,
3'h0,
3'h7,
3'h0,
3'h0,
3'h7,
3'h7,
3'h0,
3'h0,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h5,
3'h5,
3'h7,
3'h7,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h2,
3'h2,
3'h3,
3'h2,
3'h2,
3'h2,
3'h7,
3'h7,
3'h7,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h7,
3'h7,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h0,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h0,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h0,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h0,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h2,
3'h2,
3'h2,
3'h2,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h3,
3'h5,
3'h5,
3'h7,
3'h7,
3'h0,
3'h0,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h0,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h7,
3'h7,
3'h7,
3'h5,
3'h5,
3'h7,
3'h7,
3'h7,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h2,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h7,
3'h7,
3'h0,
3'h7,
3'h7,
3'h0,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h0,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h0,
3'h7,
3'h7,
3'h7,
3'h0,
3'h0,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h0,
3'h0,
3'h0,
3'h0,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h0,
3'h7,
3'h7,
3'h0,
3'h0,
3'h7,
3'h7,
3'h0,
3'h0,
3'h0,
3'h7,
3'h7,
3'h7,
3'h3,
3'h2,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h2,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h2,
3'h2,
3'h2,
3'h2,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h7,
3'h7,
3'h0,
3'h0,
3'h7,
3'h7,
3'h7,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h0,
3'h7,
3'h0,
3'h0,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h0,
3'h7,
3'h7,
3'h7,
3'h0,
3'h0,
3'h0,
3'h0,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h0,
3'h0,
3'h7,
3'h7,
3'h0,
3'h7,
3'h0,
3'h0,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h0,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h0,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h0,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h0,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h0,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h0,
3'h7,
3'h7,
3'h0,
3'h7,
3'h0,
3'h0,
3'h7,
3'h7,
3'h0,
3'h0,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h3,
3'h3,
3'h3,
3'h7,
3'h5,
3'h5,
3'h7,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h3,
3'h7,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h7,
3'h7,
3'h7,
3'h5,
3'h5,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h0,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h0,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h0,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h0,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h0,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h3,
3'h3,
3'h2,
3'h2,
3'h3,
3'h3,
3'h3,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h2,
3'h2,
3'h3,
3'h2,
3'h2,
3'h2,
3'h2,
3'h3,
3'h2,
3'h2,
3'h5,
3'h0,
3'h0,
3'h0,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h0,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h7,
3'h7,
3'h7,
3'h7,
3'h5,
3'h7,
3'h5,
3'h7,
3'h7,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h2,
3'h2,
3'h3,
3'h2,
3'h2,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h2,
3'h7,
3'h5,
3'h5,
3'h7,
3'h7,
3'h0,
3'h0,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h0,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h0,
3'h7,
3'h7,
3'h7,
3'h7,
3'h0,
3'h7,
3'h7,
3'h7,
3'h7,
3'h0,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h5,
3'h5,
3'h5,
3'h7,
3'h7,
3'h7,
3'h0,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h0,
3'h7,
3'h0,
3'h7,
3'h7,
3'h0,
3'h0,
3'h7,
3'h7,
3'h7,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h7,
3'h3,
3'h3,
3'h2,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h2,
3'h2,
3'h2,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h5,
3'h3,
3'h3,
3'h3,
3'h5,
3'h5,
3'h5,
3'h7,
3'h7,
3'h7,
3'h0,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h7,
3'h7,
3'h7,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h0,
3'h0,
3'h7,
3'h7,
3'h0,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h0,
3'h7,
3'h7,
3'h7,
3'h0,
3'h7,
3'h0,
3'h0,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h0,
3'h0,
3'h7,
3'h7,
3'h0,
3'h7,
3'h0,
3'h5,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h0,
3'h0,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h0,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h0,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h0,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h0,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h0,
3'h7,
3'h0,
3'h0,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h3,
3'h3,
3'h3,
3'h3,
3'h7,
3'h7,
3'h3,
3'h3,
3'h3,
3'h3,
3'h2,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h2,
3'h2,
3'h2,
3'h2,
3'h3,
3'h3,
3'h3,
3'h2,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h5,
3'h5,
3'h7,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h0,
3'h0,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h0,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h0,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h3,
3'h7,
3'h5,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h5,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h0,
3'h7,
3'h7,
3'h0,
3'h7,
3'h7,
3'h0,
3'h7,
3'h7,
3'h7,
3'h7,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h2,
3'h2,
3'h2,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h5,
3'h5,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h3,
3'h2,
3'h3,
3'h3,
3'h3,
3'h5,
3'h5,
3'h7,
3'h7,
3'h7,
3'h0,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h7,
3'h0,
3'h0,
3'h7,
3'h7,
3'h0,
3'h7,
3'h7,
3'h0,
3'h7,
3'h0,
3'h0,
3'h7,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h2,
3'h2,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h7,
3'h7,
3'h7,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h7,
3'h7,
3'h7,
3'h0,
3'h0,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h7,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h7,
3'h3,
3'h3,
3'h7,
3'h7,
3'h7,
3'h5,
3'h7,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h0,
3'h0,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h0,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h0,
3'h7,
3'h0,
3'h0,
3'h0,
3'h7,
3'h0,
3'h7,
3'h7,
3'h7,
3'h5,
3'h5,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h0,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h0,
3'h7,
3'h7,
3'h7,
3'h7,
3'h0,
3'h0,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h2,
3'h2,
3'h2,
3'h3,
3'h3,
3'h3,
3'h2,
3'h2,
3'h3,
3'h3,
3'h3,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h0,
3'h0,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h3,
3'h3,
3'h7,
3'h7,
3'h7,
3'h0,
3'h0,
3'h0,
3'h7,
3'h7,
3'h5,
3'h5,
3'h7,
3'h3,
3'h3,
3'h3,
3'h3,
3'h7,
3'h5,
3'h5,
3'h7,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h7,
3'h7,
3'h7,
3'h0,
3'h5,
3'h7,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h7,
3'h5,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h0,
3'h7,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h2,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h7,
3'h0,
3'h0,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h0,
3'h7,
3'h7,
3'h5,
3'h7,
3'h7,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h7,
3'h5,
3'h7,
3'h3,
3'h3,
3'h7,
3'h5,
3'h5,
3'h7,
3'h7,
3'h3,
3'h3,
3'h3,
3'h3,
3'h7,
3'h7,
3'h0,
3'h0,
3'h0,
3'h0,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h5,
3'h5,
3'h7,
3'h3,
3'h3,
3'h3,
3'h3,
3'h7,
3'h7,
3'h5,
3'h7,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h7,
3'h7,
3'h7,
3'h7,
3'h5,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h0,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h0,
3'h0,
3'h0,
3'h0,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h7,
3'h5,
3'h7,
3'h7,
3'h7,
3'h7,
3'h3,
3'h7,
3'h7,
3'h7,
3'h7,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h0,
3'h7,
3'h7,
3'h7,
3'h7,
3'h0,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h2,
3'h2,
3'h2,
3'h3,
3'h5,
3'h7,
3'h7,
3'h7,
3'h7,
3'h0,
3'h0,
3'h7,
3'h7,
3'h0,
3'h0,
3'h0,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h0,
3'h0,
3'h0,
3'h0,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h2,
3'h2,
3'h2,
3'h2,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h3,
3'h7,
3'h7,
3'h7,
3'h0,
3'h0,
3'h7,
3'h7,
3'h7,
3'h5,
3'h3,
3'h3,
3'h2,
3'h2,
3'h2,
3'h3,
3'h7,
3'h7,
3'h7,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h7,
3'h7,
3'h7,
3'h0,
3'h0,
3'h7,
3'h7,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h2,
3'h2,
3'h2,
3'h3,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h7,
3'h7,
3'h7,
3'h0,
3'h7,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h7,
3'h7,
3'h0,
3'h0,
3'h7,
3'h7,
3'h7,
3'h7,
3'h5,
3'h7,
3'h7,
3'h5,
3'h5,
3'h5,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h7,
3'h5,
3'h7,
3'h7,
3'h7,
3'h7,
3'h5,
3'h5,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h0,
3'h0,
3'h0,
3'h0,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h5,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h0,
3'h0,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h0,
3'h7,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h7,
3'h7,
3'h3,
3'h3,
3'h3,
3'h3,
3'h2,
3'h3,
3'h7,
3'h7,
3'h7,
3'h7,
3'h0,
3'h0,
3'h0,
3'h0,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h7,
3'h7,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h2,
3'h2,
3'h3,
3'h5,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h0,
3'h0,
3'h0,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h5,
3'h5,
3'h7,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h3,
3'h3,
3'h3,
3'h3,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h3,
3'h3,
3'h3,
3'h7,
3'h7,
3'h7,
3'h0,
3'h7,
3'h7,
3'h3,
3'h3,
3'h3,
3'h3,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h7,
3'h7,
3'h0,
3'h0,
3'h0,
3'h0,
3'h7,
3'h7,
3'h0,
3'h7,
3'h7,
3'h7,
3'h5,
3'h7,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h7,
3'h3,
3'h3,
3'h3,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h5,
3'h7,
3'h3,
3'h2,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h7,
3'h7,
3'h7,
3'h7,
3'h0,
3'h7,
3'h7,
3'h7,
3'h7,
3'h0,
3'h0,
3'h7,
3'h7,
3'h7,
3'h0,
3'h7,
3'h7,
3'h5,
3'h7,
3'h7,
3'h7,
3'h3,
3'h7,
3'h7,
3'h7,
3'h5,
3'h5,
3'h5,
3'h5,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h5,
3'h7,
3'h7,
3'h7,
3'h7,
3'h5,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h7,
3'h7,
3'h7,
3'h0,
3'h0,
3'h0,
3'h0,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h5,
3'h5,
3'h7,
3'h7,
3'h7,
3'h5,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h0,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h0,
3'h7,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h0,
3'h7,
3'h0,
3'h0,
3'h7,
3'h7,
3'h7,
3'h7,
3'h3,
3'h3,
3'h3,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h3,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h3,
3'h3,
3'h5,
3'h7,
3'h7,
3'h7,
3'h7,
3'h0,
3'h0,
3'h0,
3'h0,
3'h7,
3'h0,
3'h7,
3'h7,
3'h7,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h7,
3'h7,
3'h7,
3'h7,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h0,
3'h0,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h0,
3'h0,
3'h0,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h2,
3'h3,
3'h2,
3'h2,
3'h3,
3'h3,
3'h3,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h7,
3'h7,
3'h7,
3'h7,
3'h3,
3'h3,
3'h3,
3'h3,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h7,
3'h5,
3'h0,
3'h7,
3'h0,
3'h0,
3'h7,
3'h7,
3'h0,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h2,
3'h2,
3'h2,
3'h2,
3'h3,
3'h3,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h0,
3'h0,
3'h0,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h5,
3'h0,
3'h0,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h0,
3'h7,
3'h7,
3'h7,
3'h7,
3'h3,
3'h2,
3'h2,
3'h2,
3'h2,
3'h7,
3'h5,
3'h7,
3'h5,
3'h7,
3'h7,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h7,
3'h7,
3'h5,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h7,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h0,
3'h7,
3'h0,
3'h5,
3'h7,
3'h7,
3'h7,
3'h3,
3'h3,
3'h3,
3'h3,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h3,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h0,
3'h0,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h3,
3'h3,
3'h3,
3'h3,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h0,
3'h7,
3'h7,
3'h7,
3'h7,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h0,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h2,
3'h2,
3'h2,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h3,
3'h5,
3'h5,
3'h5,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h0,
3'h7,
3'h7,
3'h3,
3'h3,
3'h3,
3'h3,
3'h7,
3'h7,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h3,
3'h5,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h0,
3'h7,
3'h7,
3'h5,
3'h7,
3'h7,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h5,
3'h7,
3'h3,
3'h3,
3'h3,
3'h3,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h3,
3'h7,
3'h5,
3'h7,
3'h7,
3'h7,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h7,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h0,
3'h0,
3'h0,
3'h0,
3'h7,
3'h7,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h0,
3'h0,
3'h7,
3'h7,
3'h0,
3'h0,
3'h0,
3'h0,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h0,
3'h0,
3'h0,
3'h0,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h3,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h3,
3'h3,
3'h3,
3'h3,
3'h2,
3'h3,
3'h3,
3'h3,
3'h3,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h0,
3'h0,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h3,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h5,
3'h7,
3'h7,
3'h7,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h7,
3'h7,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h7,
3'h7,
3'h7,
3'h7,
3'h0,
3'h0,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h0,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h2,
3'h2,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h2,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h3,
3'h3,
3'h5,
3'h5,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h0,
3'h7,
3'h7,
3'h3,
3'h3,
3'h3,
3'h3,
3'h7,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h2,
3'h2,
3'h3,
3'h3,
3'h2,
3'h2,
3'h2,
3'h5,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h0,
3'h7,
3'h7,
3'h7,
3'h0,
3'h0,
3'h0,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h3,
3'h3,
3'h3,
3'h3,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h7,
3'h5,
3'h7,
3'h7,
3'h7,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h0,
3'h0,
3'h0,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h0,
3'h0,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h0,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h0,
3'h7,
3'h0,
3'h0,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h0,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h0,
3'h0,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h0,
3'h0,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h3,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h0,
3'h0,
3'h7,
3'h7,
3'h7,
3'h3,
3'h3,
3'h3,
3'h3,
3'h7,
3'h7,
3'h7,
3'h7,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h7,
3'h7,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h5,
3'h0,
3'h7,
3'h0,
3'h0,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h2,
3'h2,
3'h2,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h5,
3'h5,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h2,
3'h2,
3'h2,
3'h3,
3'h2,
3'h2,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h0,
3'h0,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h3,
3'h3,
3'h3,
3'h2,
3'h3,
3'h3,
3'h2,
3'h3,
3'h2,
3'h2,
3'h3,
3'h3,
3'h3,
3'h5,
3'h7,
3'h7,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h0,
3'h7,
3'h0,
3'h0,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h0,
3'h0,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h0,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h0,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h0,
3'h0,
3'h7,
3'h7,
3'h7,
3'h7,
3'h0,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h0,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h0,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h0,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h0,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h2,
3'h2,
3'h2,
3'h2,
3'h3,
3'h7,
3'h7,
3'h7,
3'h7,
3'h5,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h5,
3'h5,
3'h3,
3'h2,
3'h3,
3'h3,
3'h3,
3'h3,
3'h7,
3'h5,
3'h5,
3'h7,
3'h7,
3'h7,
3'h0,
3'h0,
3'h7,
3'h7,
3'h0,
3'h0,
3'h7,
3'h7,
3'h5,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h0,
3'h0,
3'h7,
3'h5,
3'h5,
3'h7,
3'h3,
3'h3,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h7,
3'h7,
3'h7,
3'h0,
3'h0,
3'h0,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h3,
3'h3,
3'h7,
3'h7,
3'h5,
3'h0,
3'h7,
3'h7,
3'h7,
3'h7,
3'h0,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h0,
3'h7,
3'h7,
3'h0,
3'h7,
3'h7,
3'h7,
3'h7,
3'h0,
3'h5,
3'h7,
3'h7,
3'h7,
3'h7,
3'h0,
3'h7,
3'h0,
3'h0,
3'h7,
3'h7,
3'h7,
3'h0,
3'h0,
3'h0,
3'h7,
3'h0,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h0,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h7,
3'h5,
3'h5,
3'h3,
3'h3,
3'h3,
3'h2,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h2,
3'h2,
3'h2,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h2,
3'h2,
3'h2,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h0,
3'h7,
3'h0,
3'h7,
3'h7,
3'h0,
3'h7,
3'h7,
3'h7,
3'h7,
3'h0,
3'h7,
3'h7,
3'h7,
3'h7,
3'h0,
3'h7,
3'h7,
3'h0,
3'h7,
3'h7,
3'h0,
3'h7,
3'h7,
3'h7,
3'h7,
3'h0,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h5,
3'h5,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h7,
3'h5,
3'h5,
3'h7,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h7,
3'h7,
3'h7,
3'h7,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h0,
3'h7,
3'h7,
3'h0,
3'h7,
3'h7,
3'h7,
3'h7,
3'h0,
3'h7,
3'h7,
3'h0,
3'h7,
3'h0,
3'h7,
3'h7,
3'h0,
3'h7,
3'h7,
3'h0,
3'h7,
3'h0,
3'h7,
3'h7,
3'h0,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h0,
3'h7,
3'h0,
3'h7,
3'h7,
3'h0,
3'h7,
3'h0,
3'h7,
3'h7,
3'h7,
3'h0,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h0,
3'h7,
3'h7,
3'h0,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h0,
3'h0,
3'h7,
3'h0,
3'h7,
3'h7,
3'h0,
3'h7,
3'h7,
3'h7,
3'h7,
3'h0,
3'h7,
3'h7,
3'h7,
3'h7,
3'h0,
3'h0,
3'h7,
3'h7,
3'h7,
3'h7,
3'h0,
3'h7,
3'h7,
3'h7,
3'h7,
3'h0,
3'h7,
3'h7,
3'h7,
3'h7,
3'h0,
3'h0,
3'h7,
3'h0,
3'h7,
3'h7,
3'h0,
3'h7,
3'h7,
3'h7,
3'h7,
3'h0,
3'h7,
3'h7,
3'h7,
3'h7,
3'h0,
3'h0,
3'h7,
3'h0,
3'h7,
3'h7,
3'h0,
3'h7,
3'h0,
3'h7,
3'h7,
3'h7,
3'h5,
3'h7,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h2,
3'h2,
3'h2,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h5,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h0,
3'h7,
3'h7,
3'h7,
3'h0,
3'h0,
3'h7,
3'h7,
3'h7,
3'h0,
3'h0,
3'h7,
3'h0,
3'h7,
3'h7,
3'h0,
3'h7,
3'h7,
3'h7,
3'h7,
3'h0,
3'h7,
3'h7,
3'h7,
3'h7,
3'h0,
3'h0,
3'h7,
3'h0,
3'h7,
3'h7,
3'h0,
3'h7,
3'h7,
3'h7,
3'h7,
3'h0,
3'h7,
3'h7,
3'h7,
3'h7,
3'h0,
3'h7,
3'h7,
3'h0,
3'h7,
3'h7,
3'h0,
3'h7,
3'h7,
3'h0,
3'h7,
3'h0,
3'h7,
3'h7,
3'h0,
3'h7,
3'h7,
3'h7,
3'h7,
3'h0,
3'h7,
3'h7,
3'h7,
3'h7,
3'h0,
3'h0,
3'h7,
3'h0,
3'h7,
3'h7,
3'h0,
3'h7,
3'h7,
3'h7,
3'h7,
3'h0,
3'h7,
3'h7,
3'h7,
3'h7,
3'h0,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h5,
3'h7,
3'h7,
3'h7,
3'h7,
3'h5,
3'h7,
3'h7,
3'h0,
3'h7,
3'h7,
3'h0,
3'h7,
3'h0,
3'h7,
3'h7,
3'h0,
3'h7,
3'h7,
3'h7,
3'h7,
3'h0,
3'h7,
3'h7,
3'h7,
3'h7,
3'h0,
3'h0,
3'h7,
3'h7,
3'h7,
3'h7,
3'h5,
3'h7,
3'h7,
3'h7,
3'h7,
3'h0,
3'h7,
3'h7,
3'h7,
3'h3,
3'h7,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h7,
3'h3,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h0,
3'h7,
3'h7,
3'h0,
3'h7,
3'h7,
3'h0,
3'h7,
3'h0,
3'h7,
3'h7,
3'h0,
3'h7,
3'h7,
3'h7,
3'h7,
3'h0,
3'h7,
3'h7,
3'h7,
3'h7,
3'h0,
3'h0,
3'h7,
3'h0,
3'h7,
3'h7,
3'h0,
3'h7,
3'h7,
3'h7,
3'h7,
3'h0,
3'h7,
3'h7,
3'h7,
3'h7,
3'h0,
3'h0,
3'h7,
3'h0,
3'h7,
3'h7,
3'h0,
3'h7,
3'h7,
3'h7,
3'h7,
3'h0,
3'h7,
3'h7,
3'h0,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h3,
3'h3,
3'h3,
3'h3,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h0,
3'h7,
3'h0,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h5,
3'h7,
3'h7,
3'h7,
3'h7,
3'h0,
3'h7,
3'h7,
3'h7,
3'h0,
3'h0,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h7,
3'h7,
3'h7,
3'h5,
3'h7,
3'h7,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h2,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h2,
3'h2,
3'h3,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h7,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h2,
3'h2,
3'h3,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h0,
3'h7,
3'h7,
3'h7,
3'h7,
3'h0,
3'h7,
3'h7,
3'h7,
3'h7,
3'h0,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h0,
3'h7,
3'h7,
3'h7,
3'h7,
3'h0,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h3,
3'h3,
3'h3,
3'h3,
3'h5,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h3,
3'h5,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h0,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h0,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h0,
3'h7,
3'h7,
3'h7,
3'h7,
3'h0,
3'h7,
3'h7,
3'h0,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h0,
3'h7,
3'h7,
3'h7,
3'h7,
3'h0,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h0,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h0,
3'h7,
3'h7,
3'h7,
3'h7,
3'h0,
3'h7,
3'h7,
3'h7,
3'h7,
3'h0,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h0,
3'h7,
3'h7,
3'h7,
3'h7,
3'h0,
3'h7,
3'h7,
3'h7,
3'h7,
3'h0,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h0,
3'h7,
3'h7,
3'h7,
3'h7,
3'h0,
3'h7,
3'h7,
3'h7,
3'h7,
3'h0,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h0,
3'h7,
3'h7,
3'h7,
3'h7,
3'h0,
3'h7,
3'h7,
3'h7,
3'h7,
3'h5,
3'h7,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h2,
3'h2,
3'h3,
3'h3,
3'h3,
3'h3,
3'h2,
3'h2,
3'h3,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h0,
3'h0,
3'h7,
3'h0,
3'h7,
3'h0,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h0,
3'h7,
3'h7,
3'h7,
3'h7,
3'h0,
3'h7,
3'h7,
3'h7,
3'h7,
3'h0,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h0,
3'h7,
3'h7,
3'h7,
3'h7,
3'h0,
3'h7,
3'h7,
3'h7,
3'h7,
3'h0,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h0,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h0,
3'h7,
3'h7,
3'h7,
3'h7,
3'h0,
3'h7,
3'h7,
3'h7,
3'h7,
3'h0,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h0,
3'h7,
3'h7,
3'h7,
3'h7,
3'h0,
3'h7,
3'h7,
3'h7,
3'h7,
3'h0,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h0,
3'h7,
3'h7,
3'h7,
3'h7,
3'h0,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h0,
3'h7,
3'h7,
3'h7,
3'h7,
3'h0,
3'h7,
3'h7,
3'h7,
3'h7,
3'h0,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h0,
3'h7,
3'h7,
3'h7,
3'h7,
3'h0,
3'h7,
3'h7,
3'h0,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h0,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h0,
3'h7,
3'h7,
3'h7,
3'h7,
3'h0,
3'h7,
3'h7,
3'h7,
3'h7,
3'h0,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h0,
3'h7,
3'h7,
3'h7,
3'h7,
3'h0,
3'h7,
3'h7,
3'h7,
3'h7,
3'h0,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h0,
3'h7,
3'h7,
3'h7,
3'h7,
3'h0,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h0,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h3,
3'h3,
3'h3,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h2,
3'h2,
3'h3,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h3,
3'h3,
3'h3,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h3,
3'h3,
3'h3,
3'h3,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h2,
3'h2,
3'h3,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h0,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h2,
3'h2,
3'h2,
3'h3,
3'h3,
3'h3,
3'h3,
3'h2,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h3,
3'h3,
3'h3,
3'h3,
3'h7,
3'h7,
3'h7,
3'h3,
3'h7,
3'h3,
3'h5,
3'h7,
3'h7,
3'h0,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h0,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h0,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h0,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h0,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h0,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h2,
3'h2,
3'h2,
3'h3,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h0,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h0,
3'h7,
3'h7,
3'h7,
3'h7,
3'h0,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h0,
3'h7,
3'h7,
3'h0,
3'h7,
3'h7,
3'h7,
3'h7,
3'h5,
3'h7,
3'h7,
3'h7,
3'h7,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h7,
3'h5,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h2,
3'h2,
3'h3,
3'h3,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h2,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h2,
3'h2,
3'h3,
3'h3,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h5,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h0,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h0,
3'h7,
3'h7,
3'h0,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h2,
3'h2,
3'h3,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h0,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h5,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h7,
3'h5,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h0,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h3,
3'h3,
3'h3,
3'h7,
3'h7,
3'h7,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h7,
3'h7,
3'h7,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h7,
3'h7,
3'h7,
3'h7,
3'h5,
3'h7,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h0,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h7,
3'h7,
3'h5,
3'h5,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h0,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h2,
3'h2,
3'h2,
3'h3,
3'h5,
3'h5,
3'h5,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h5,
3'h5,
3'h7,
3'h5,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h0,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h0,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h3,
3'h3,
3'h3,
3'h5,
3'h7,
3'h5,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h5,
3'h7,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h5,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h0,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h0,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h5,
3'h7,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h7,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h0,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h5,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h7,
3'h7,
3'h7,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h0,
3'h7,
3'h7,
3'h7,
3'h7,
3'h0,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h2,
3'h3,
3'h3,
3'h3,
3'h3,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h0,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h0,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h5,
3'h7,
3'h7,
3'h3,
3'h3,
3'h3,
3'h3,
3'h7,
3'h7,
3'h7,
3'h7,
3'h5,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h5,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h5,
3'h7,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h5,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h0,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h0,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h0,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h5,
3'h5,
3'h7,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h7,
3'h5,
3'h5,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h7,
3'h7,
3'h7,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h7,
3'h7,
3'h7,
3'h3,
3'h7,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h3,
3'h3,
3'h3,
3'h7,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h7,
3'h5,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h7,
3'h7,
3'h7,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h2,
3'h3,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h0,
3'h7,
3'h0,
3'h7,
3'h7,
3'h0,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h0,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h0,
3'h7,
3'h7,
3'h7,
3'h7,
3'h0,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h5,
3'h7,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h2,
3'h3,
3'h3,
3'h7,
3'h5,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h5,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h3,
3'h3,
3'h7,
3'h3,
3'h3,
3'h3,
3'h3,
3'h7,
3'h7,
3'h3,
3'h7,
3'h7,
3'h7,
3'h3,
3'h7,
3'h7,
3'h5,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h5,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h0,
3'h7,
3'h7,
3'h7,
3'h7,
3'h0,
3'h7,
3'h7,
3'h0,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h0,
3'h7,
3'h7,
3'h0,
3'h7,
3'h7,
3'h7,
3'h7,
3'h0,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h5,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h7,
3'h7,
3'h7,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h3,
3'h3,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h7,
3'h7,
3'h5,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h3,
3'h3,
3'h7,
3'h5,
3'h7,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h2,
3'h3,
3'h3,
3'h3,
3'h3,
3'h7,
3'h7,
3'h5,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h5,
3'h7,
3'h7,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h7,
3'h3,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h2,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h0,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h0,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h0,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h5,
3'h7,
3'h7,
3'h0,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h5,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h3,
3'h3,
3'h3,
3'h7,
3'h7,
3'h7,
3'h7,
3'h3,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h5,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h0,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h3,
3'h3,
3'h3,
3'h3,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h0,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h5,
3'h3,
3'h3,
3'h3,
3'h3,
3'h7,
3'h3,
3'h3,
3'h3,
3'h7,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h5,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h5,
3'h5,
3'h7,
3'h3,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h3,
3'h3,
3'h3,
3'h7,
3'h7,
3'h7,
3'h7,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h5,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h7,
3'h3,
3'h7,
3'h3,
3'h7,
3'h5,
3'h7,
3'h5,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h3,
3'h3,
3'h3,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h7,
3'h5,
3'h5,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h5,
3'h7,
3'h3,
3'h3,
3'h3,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h2,
3'h5,
3'h7,
3'h7,
3'h7,
3'h7,
3'h5,
3'h5,
3'h5,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h5,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h5,
3'h7,
3'h7,
3'h5,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h0,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h5,
3'h7,
3'h3,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h0,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h3,
3'h5,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h5,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h7,
3'h5,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h3,
3'h3,
3'h2,
3'h3,
3'h3,
3'h3,
3'h3,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h3,
3'h3,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h5,
3'h7,
3'h7,
3'h5,
3'h7,
3'h7,
3'h5,
3'h7,
3'h5,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h3,
3'h3,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h5,
3'h7,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h5,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h5,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h3,
3'h3,
3'h3,
3'h3,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h3,
3'h2,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h3,
3'h3,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h3,
3'h3,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h3,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h3,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h3,
3'h3,
3'h2,
3'h2,
3'h2,
3'h2,
3'h3,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h3,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h3,
3'h2,
3'h3,
3'h3,
3'h2,
3'h2,
3'h2,
3'h3,
3'h3,
3'h3,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h3,
3'h2,
3'h2,
3'h2,
3'h3,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h3,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h3,
3'h2,
3'h2,
3'h2,
3'h3,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h3,
3'h3,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h3,
3'h2,
3'h2,
3'h3,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h3,
3'h3,
3'h2,
3'h3,
3'h3,
3'h2,
3'h2,
3'h3,
3'h2,
3'h2,
3'h2,
3'h3,
3'h3,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h3,
3'h2,
3'h2,
3'h2,
3'h3,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h3,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h3,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h3,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h3,
3'h3,
3'h2,
3'h2,
3'h3,
3'h3,
3'h2,
3'h2,
3'h3,
3'h3,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h3,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h3,
3'h2,
3'h3,
3'h3,
3'h2,
3'h2,
3'h3,
3'h3,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h3,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h3,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h3,
3'h3,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h3,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h3,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h3,
3'h3,
3'h2,
3'h2,
3'h2,
3'h2,
3'h3,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h3,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h3,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h3,
3'h3,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h3,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h3,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h3,
3'h3,
3'h2,
3'h2,
3'h2,
3'h2,
3'h3,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h3,
3'h2,
3'h3,
3'h2,
3'h2,
3'h3,
3'h2,
3'h2,
3'h2,
3'h2,
3'h3,
3'h3,
3'h2,
3'h3,
3'h2,
3'h2,
3'h2,
3'h2,
3'h3,
3'h3,
3'h2,
3'h2,
3'h2,
3'h3,
3'h3,
3'h2,
3'h2,
3'h2,
3'h2,
3'h3,
3'h3,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h3,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h3,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h3,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h3,
3'h3,
3'h2,
3'h2,
3'h2,
3'h2,
3'h3,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h2,
3'h3,
3'h2,
3'h2,
3'h2,
3'h3,
3'h2,
3'h2,
3'h5,
3'h5,
3'h5,
3'h3,
3'h3,
3'h5,
3'h5,
3'h3,
3'h2,
3'h3,
3'h5,
3'h5,
3'h5,
3'h5,
3'h5,
3'h5,
3'h5,
3'h5,
3'h3,
3'h3,
3'h5,
3'h5,
3'h5,
3'h5,
3'h5,
3'h5,
3'h5,
3'h3,
3'h3,
3'h3,
3'h5,
3'h5,
3'h3,
3'h3,
3'h5,
3'h5,
3'h5,
3'h5,
3'h5,
3'h3,
3'h3,
3'h5,
3'h5,
3'h5,
3'h5,
3'h5,
3'h5,
3'h3,
3'h3,
3'h5,
3'h5,
3'h5,
3'h5,
3'h5,
3'h5,
3'h5,
3'h5,
3'h5,
3'h3,
3'h3,
3'h5,
3'h5,
3'h5,
3'h5,
3'h5,
3'h5,
3'h5,
3'h3,
3'h3,
3'h3,
3'h5,
3'h5,
3'h5,
3'h3,
3'h5,
3'h5,
3'h5,
3'h5,
3'h3,
3'h5,
3'h3,
3'h3,
3'h3,
3'h5,
3'h5,
3'h5,
3'h5,
3'h5,
3'h5,
3'h5,
3'h3,
3'h3,
3'h5,
3'h5,
3'h5,
3'h3,
3'h5,
3'h5,
3'h5,
3'h5,
3'h5,
3'h3,
3'h3,
3'h5,
3'h3,
3'h5,
3'h5,
3'h5,
3'h5,
3'h3,
3'h3,
3'h5,
3'h5,
3'h5,
3'h5,
3'h5,
3'h3,
3'h3,
3'h5,
3'h5,
3'h3,
3'h3,
3'h3,
3'h5,
3'h5,
3'h5,
3'h5,
3'h5,
3'h5,
3'h5,
3'h3,
3'h3,
3'h5,
3'h5,
3'h5,
3'h5,
3'h5,
3'h5,
3'h5,
3'h5,
3'h5,
3'h3,
3'h3,
3'h5,
3'h5,
3'h7,
3'h3,
3'h7,
3'h5,
3'h5,
3'h5,
3'h3,
3'h3,
3'h3,
3'h5,
3'h5,
3'h5,
3'h5,
3'h3,
3'h5,
3'h5,
3'h5,
3'h3,
3'h3,
3'h3,
3'h3,
3'h5,
3'h5,
3'h5,
3'h3,
3'h5,
3'h5,
3'h5,
3'h3,
3'h5,
3'h3,
3'h5,
3'h5,
3'h3,
3'h5,
3'h5,
3'h5,
3'h5,
3'h3,
3'h3,
3'h5,
3'h5,
3'h5,
3'h3,
3'h3,
3'h3,
3'h5,
3'h5,
3'h3,
3'h3,
3'h3,
3'h5,
3'h5,
3'h5,
3'h5,
3'h5,
3'h5,
3'h3,
3'h3,
3'h5,
3'h5,
3'h3,
3'h5,
3'h3,
3'h3,
3'h3,
3'h5,
3'h5,
3'h5,
3'h5,
3'h5,
3'h3,
3'h3,
3'h5,
3'h5,
3'h3,
3'h5,
3'h5,
3'h5,
3'h5,
3'h5,
3'h5,
3'h5,
3'h5,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h3,
3'h5,
3'h3,
3'h5,
3'h5,
3'h5,
3'h5,
3'h5,
3'h3,
3'h3,
3'h5,
3'h5,
3'h3,
3'h3,
3'h5,
3'h5,
3'h5,
3'h5,
3'h5,
3'h3,
3'h5,
3'h5,
3'h3,
3'h5,
3'h5,
3'h5,
3'h5,
3'h5,
3'h5,
3'h5,
3'h5,
3'h5,
3'h5,
3'h5,
3'h3,
3'h5,
3'h5,
3'h5,
3'h3,
3'h3,
3'h5,
3'h5,
3'h5,
3'h3,
3'h3,
3'h5,
3'h5,
3'h5,
3'h5,
3'h5,
3'h3,
3'h5,
3'h5,
3'h3,
3'h3,
3'h3,
3'h3,
3'h5,
3'h5,
3'h3,
3'h3,
3'h5,
3'h5,
3'h3,
3'h3,
3'h3,
3'h3,
3'h5,
3'h5,
3'h5,
3'h3,
3'h5,
3'h3,
3'h3,
3'h5,
3'h5,
3'h3,
3'h3,
3'h5,
3'h5,
3'h5,
3'h5,
3'h3,
3'h3,
3'h5,
3'h5,
3'h3,
3'h2,
3'h3,
3'h5,
3'h5,
3'h5,
3'h5,
3'h5,
3'h5,
3'h5,
3'h5,
3'h3,
3'h3,
3'h5,
3'h5,
3'h5,
3'h5,
3'h5,
3'h5,
3'h5,
3'h3,
3'h3,
3'h3,
3'h5,
3'h5,
3'h3,
3'h3,
3'h5,
3'h5,
3'h5,
3'h5,
3'h5,
3'h3,
3'h3,
3'h5,
3'h5,
3'h5,
3'h5,
3'h5,
3'h5,
3'h3,
3'h3,
3'h5,
3'h5,
3'h5,
3'h5,
3'h5,
3'h5,
3'h5,
3'h5,
3'h5,
3'h3,
3'h3,
3'h5,
3'h5,
3'h5,
3'h5,
3'h5,
3'h5,
3'h5,
3'h3,
3'h3,
3'h3,
3'h5,
3'h5,
3'h3,
3'h5,
3'h5,
3'h5,
3'h5,
3'h5,
3'h3,
3'h3,
3'h3,
3'h5,
3'h5,
3'h3,
3'h3,
3'h5,
3'h5,
3'h5,
3'h5,
3'h5,
3'h5,
3'h5,
3'h3,
3'h3,
3'h3,
3'h5,
3'h5,
3'h5,
3'h5,
3'h5,
3'h5,
3'h5,
3'h5,
3'h3,
3'h5,
3'h3,
3'h3,
3'h5,
3'h5,
3'h3,
3'h3,
3'h5,
3'h5,
3'h5,
3'h5,
3'h3,
3'h3,
3'h5,
3'h5,
3'h3,
3'h2,
3'h3,
3'h5,
3'h5,
3'h5,
3'h5,
3'h5,
3'h5,
3'h5,
3'h5,
3'h3,
3'h3,
3'h5,
3'h5,
3'h5,
3'h5,
3'h5,
3'h5,
3'h5,
3'h3,
3'h3,
3'h3,
3'h5,
3'h5,
3'h3,
3'h3,
3'h5,
3'h5,
3'h5,
3'h5,
3'h5,
3'h3,
3'h3,
3'h5,
3'h5,
3'h5,
3'h5,
3'h5,
3'h5,
3'h3,
3'h3,
3'h5,
3'h5,
3'h5,
3'h5,
3'h5,
3'h5,
3'h5,
3'h5,
3'h5,
3'h3,
3'h3,
3'h5,
3'h5,
3'h5,
3'h5,
3'h5,
3'h5,
3'h5,
3'h3,
3'h3,
3'h3,
3'h5,
3'h5,
3'h3,
3'h3,
3'h5,
3'h5,
3'h5,
3'h5,
3'h5,
3'h5,
3'h5,
3'h5,
3'h5,
3'h5,
3'h5,
3'h3,
3'h3,
3'h5,
3'h5,
3'h5,
3'h5,
3'h5,
3'h5,
3'h5,
3'h3,
3'h3,
3'h5,
3'h5,
3'h5,
3'h3,
3'h5,
3'h5,
3'h5,
3'h5,
3'h5,
3'h5,
3'h3,
3'h3,
3'h5,
3'h5,
3'h5,
3'h3,
3'h5,
3'h5,
3'h3,
3'h3,
3'h5,
3'h5,
3'h5,
3'h5,
3'h3,
3'h5,
3'h5,
3'h5,
3'h5,
3'h3,
3'h3,
3'h5,
3'h5,
3'h5,
3'h5,
3'h5,
3'h5,
3'h3,
3'h3,
3'h3,
3'h3,
3'h5,
3'h5,
3'h5,
3'h5,
3'h5,
3'h5,
3'h5,
3'h5,
3'h5,
3'h3,
3'h3,
3'h5,
3'h5,
3'h5,
3'h5,
3'h5,
3'h5,
3'h5,
3'h3,
3'h3,
3'h3,
3'h5,
3'h5,
3'h3,
3'h3,
3'h5,
3'h5,
3'h5,
3'h5,
3'h5,
3'h3,
3'h3,
3'h5,
3'h5,
3'h5,
3'h5,
3'h5,
3'h5,
3'h3,
3'h3,
3'h5,
3'h5,
3'h5,
3'h5,
3'h5,
3'h5,
3'h5,
3'h5,
3'h5,
3'h3,
3'h3,
3'h5,
3'h5,
3'h5,
3'h5,
3'h5,
3'h5,
3'h5,
3'h3,
3'h3,
3'h3,
3'h5,
3'h5,
3'h5,
3'h5,
3'h5,
3'h3,
3'h5,
3'h5,
3'h5,
3'h5,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h5,
3'h7,
3'h7,
3'h7,
3'h7,
3'h5,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h5,
3'h5,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h5,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h5,
3'h7,
3'h7,
3'h7,
3'h5,
3'h7,
3'h7,
3'h7,
3'h7,
3'h5,
3'h5,
3'h7,
3'h7,
3'h7,
3'h5,
3'h5,
3'h7,
3'h7,
3'h7,
3'h5,
3'h7,
3'h7,
3'h5,
3'h5,
3'h7,
3'h7,
3'h7,
3'h5,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h5,
3'h5,
3'h5,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h5,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h5,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h5,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h5,
3'h7,
3'h7,
3'h7,
3'h7,
3'h5,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h5,
3'h5,
3'h7,
3'h7,
3'h5,
3'h5,
3'h5,
3'h5,
3'h5,
3'h5,
3'h7,
3'h7,
3'h5,
3'h5,
3'h5,
3'h5,
3'h5,
3'h7,
3'h7,
3'h5,
3'h5,
3'h5,
3'h5,
3'h5,
3'h5,
3'h5,
3'h5,
3'h5,
3'h5,
3'h5,
3'h5,
3'h5,
3'h5,
3'h5,
3'h5,
3'h5,
3'h5,
3'h5,
3'h5,
3'h5,
3'h5,
3'h5,
3'h5,
3'h5,
3'h5,
3'h5,
3'h5,
3'h5,
3'h5,
3'h5,
3'h5,
3'h5,
3'h5,
3'h5,
3'h5,
3'h5,
3'h5,
3'h5,
3'h5,
3'h5,
3'h5,
3'h3,
3'h3,
3'h5,
3'h5,
3'h5,
3'h5,
3'h5,
3'h7,
3'h5,
3'h5,
3'h5,
3'h5,
3'h5,
3'h5,
3'h7,
3'h5,
3'h5,
3'h5,
3'h5,
3'h5,
3'h7,
3'h7,
3'h7,
3'h7,
3'h5,
3'h5,
3'h7,
3'h7,
3'h7,
3'h5,
3'h7,
3'h7,
3'h7,
3'h7,
3'h5,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h5,
3'h5,
3'h7,
3'h7,
3'h5,
3'h5,
3'h7,
3'h7,
3'h7,
3'h7,
3'h5,
3'h5,
3'h5,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h5,
3'h7,
3'h7,
3'h7,
3'h7,
3'h5,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h5,
3'h5,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h5,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h5,
3'h7,
3'h7,
3'h7,
3'h5,
3'h5,
3'h7,
3'h7,
3'h7,
3'h7,
3'h5,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h5,
3'h5,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h5,
3'h7,
3'h7,
3'h7,
3'h7,
3'h5,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h5,
3'h5,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h5,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h5,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h5,
3'h7,
3'h7,
3'h7,
3'h7,
3'h5,
3'h5,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h5,
3'h5,
3'h7,
3'h7,
3'h5,
3'h5,
3'h7,
3'h7,
3'h7,
3'h5,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h5,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h5,
3'h7,
3'h7,
3'h7,
3'h7,
3'h5,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h5,
3'h5,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h5,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h7,
3'h7,
3'h7,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h7,
3'h7,
3'h0,
3'h7,
3'h7,
3'h7,
3'h0,
3'h0,
3'h0,
3'h7,
3'h0,
3'h0,
3'h0,
3'h7,
3'h7,
3'h7,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h7,
3'h7,
3'h7,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h7,
3'h7,
3'h7,
3'h7,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h7,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h7,
3'h7,
3'h7,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h7,
3'h7,
3'h0,
3'h0,
3'h7,
3'h7,
3'h7,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h7,
3'h7,
3'h7,
3'h0,
3'h0,
3'h0,
3'h0,
3'h7,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h7,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h5,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h5,
3'h5,
3'h7,
3'h7,
3'h5,
3'h5,
3'h5,
3'h5,
3'h5,
3'h5,
3'h5,
3'h5,
3'h5,
3'h5,
3'h5,
3'h5,
3'h5,
3'h5,
3'h5,
3'h5,
3'h5,
3'h5,
3'h5,
3'h5,
3'h5,
3'h5,
3'h5,
3'h5,
3'h5,
3'h5,
3'h5,
3'h5,
3'h5,
3'h5,
3'h5,
3'h5,
3'h5,
3'h5,
3'h5,
3'h5,
3'h5,
3'h5,
3'h5,
3'h5,
3'h5,
3'h5,
3'h5,
3'h5,
3'h5,
3'h5,
3'h5,
3'h5,
3'h5,
3'h5,
3'h5,
3'h5,
3'h5,
3'h5,
3'h5,
3'h5,
3'h5,
3'h5,
3'h5,
3'h5,
3'h5,
3'h5,
3'h5,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h7,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h7,
3'h7,
3'h7,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h7,
3'h7,
3'h0,
3'h7,
3'h7,
3'h7,
3'h0,
3'h0,
3'h0,
3'h7,
3'h0,
3'h0,
3'h0,
3'h7,
3'h7,
3'h7,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h7,
3'h7,
3'h7,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h7,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h7,
3'h7,
3'h0,
3'h7,
3'h7,
3'h7,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h7,
3'h7,
3'h7,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h7,
3'h7,
3'h7,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h7,
3'h7,
3'h0,
3'h7,
3'h7,
3'h7,
3'h0,
3'h0,
3'h0,
3'h7,
3'h0,
3'h0,
3'h0,
3'h7,
3'h7,
3'h7,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h7,
3'h7,
3'h7,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h7,
3'h7,
3'h7,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h7,
3'h7,
3'h7,
3'h7,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h7,
3'h7,
3'h7,
3'h7,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h7,
3'h7,
3'h7,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h7,
3'h7,
3'h0,
3'h7,
3'h7,
3'h7,
3'h0,
3'h0,
3'h0,
3'h7,
3'h0,
3'h0,
3'h0,
3'h7,
3'h7,
3'h7,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h7,
3'h7,
3'h7,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h7,
3'h7,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h7,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h7,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h7,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h7,
3'h7,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h7,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h7,
3'h7,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h7,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h7,
3'h0,
3'h0,
3'h7,
3'h7,
3'h7,
3'h7,
3'h0,
3'h0,
3'h7,
3'h0,
3'h0,
3'h0,
3'h7,
3'h7,
3'h0,
3'h0,
3'h0,
3'h0,
3'h7,
3'h7,
3'h0,
3'h0,
3'h0,
3'h7,
3'h0,
3'h0,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h5,
3'h5,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h5,
3'h7,
3'h7,
3'h5,
3'h5,
3'h5,
3'h5,
3'h5,
3'h5,
3'h5,
3'h5,
3'h5,
3'h5,
3'h5,
3'h5,
3'h5,
3'h5,
3'h5,
3'h5,
3'h5,
3'h5,
3'h5,
3'h5,
3'h5,
3'h5,
3'h5,
3'h5,
3'h5,
3'h5,
3'h5,
3'h5,
3'h5,
3'h5,
3'h5,
3'h5,
3'h5,
3'h5,
3'h5,
3'h5,
3'h5,
3'h5,
3'h5,
3'h5,
3'h5,
3'h5,
3'h5,
3'h5,
3'h5,
3'h5,
3'h5,
3'h5,
3'h5,
3'h5,
3'h5,
3'h5,
3'h7,
3'h5,
3'h7,
3'h5,
3'h5,
3'h5,
3'h5,
3'h5,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h7,
3'h0,
3'h0,
3'h0,
3'h0,
3'h7,
3'h7,
3'h0,
3'h0,
3'h7,
3'h0,
3'h0,
3'h7,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h7,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h7,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h7,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h7,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h7,
3'h0,
3'h0,
3'h7,
3'h7,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h7,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h7,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h7,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h7,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h7,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h7,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h7,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h7,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h7,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h7,
3'h0,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h0,
3'h0,
3'h0,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h0,
3'h6,
3'h6,
3'h6,
3'h0,
3'h0,
3'h0,
3'h0,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h0,
3'h0,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h0,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h0,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h0,
3'h6,
3'h0,
3'h0,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h0,
3'h6,
3'h6,
3'h6,
3'h6,
3'h0,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h0,
3'h6,
3'h6,
3'h0,
3'h0,
3'h6,
3'h6,
3'h0,
3'h6,
3'h6,
3'h0,
3'h6,
3'h6,
3'h0,
3'h6,
3'h6,
3'h6,
3'h0,
3'h6,
3'h6,
3'h6,
3'h6,
3'h0,
3'h6,
3'h6,
3'h6,
3'h6,
3'h0,
3'h0,
3'h6,
3'h6,
3'h6,
3'h6,
3'h0,
3'h6,
3'h6,
3'h6,
3'h6,
3'h0,
3'h6,
3'h0,
3'h6,
3'h6,
3'h6,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h7,
3'h7,
3'h0,
3'h0,
3'h7,
3'h7,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h7,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h5,
3'h0,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h5,
3'h7,
3'h5,
3'h5,
3'h5,
3'h5,
3'h5,
3'h5,
3'h7,
3'h7,
3'h7,
3'h7,
3'h5,
3'h5,
3'h5,
3'h5,
3'h5,
3'h5,
3'h5,
3'h7,
3'h5,
3'h5,
3'h5,
3'h5,
3'h5,
3'h5,
3'h5,
3'h5,
3'h5,
3'h7,
3'h7,
3'h5,
3'h5,
3'h5,
3'h5,
3'h5,
3'h5,
3'h7,
3'h7,
3'h5,
3'h5,
3'h7,
3'h7,
3'h5,
3'h7,
3'h5,
3'h7,
3'h7,
3'h5,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h5,
3'h5,
3'h5,
3'h7,
3'h7,
3'h0,
3'h0,
3'h0,
3'h7,
3'h7,
3'h7,
3'h7,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h7,
3'h0,
3'h7,
3'h0,
3'h0,
3'h7,
3'h0,
3'h0,
3'h0,
3'h0,
3'h7,
3'h7,
3'h7,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h6,
3'h6,
3'h6,
3'h6,
3'h0,
3'h0,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h0,
3'h0,
3'h0,
3'h0,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h0,
3'h6,
3'h6,
3'h6,
3'h0,
3'h0,
3'h0,
3'h0,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h0,
3'h0,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h0,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h0,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h0,
3'h6,
3'h0,
3'h0,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h0,
3'h6,
3'h0,
3'h0,
3'h6,
3'h6,
3'h0,
3'h6,
3'h6,
3'h0,
3'h0,
3'h6,
3'h0,
3'h0,
3'h0,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h0,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h0,
3'h0,
3'h0,
3'h0,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h0,
3'h6,
3'h6,
3'h6,
3'h0,
3'h0,
3'h0,
3'h0,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h0,
3'h0,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h0,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h0,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h0,
3'h6,
3'h0,
3'h0,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h0,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h0,
3'h6,
3'h6,
3'h6,
3'h0,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h0,
3'h0,
3'h6,
3'h6,
3'h0,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h0,
3'h0,
3'h6,
3'h6,
3'h6,
3'h0,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h0,
3'h6,
3'h6,
3'h6,
3'h0,
3'h0,
3'h0,
3'h0,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h0,
3'h0,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h0,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h0,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h0,
3'h6,
3'h0,
3'h0,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h0,
3'h6,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h6,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h6,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h6,
3'h0,
3'h0,
3'h0,
3'h6,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h6,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h6,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h6,
3'h0,
3'h0,
3'h0,
3'h0,
3'h6,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h6,
3'h0,
3'h0,
3'h6,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h6,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h7,
3'h7,
3'h0,
3'h7,
3'h7,
3'h7,
3'h0,
3'h0,
3'h0,
3'h7,
3'h7,
3'h0,
3'h0,
3'h0,
3'h7,
3'h7,
3'h7,
3'h0,
3'h7,
3'h7,
3'h7,
3'h7,
3'h0,
3'h0,
3'h0,
3'h7,
3'h0,
3'h0,
3'h5,
3'h7,
3'h7,
3'h7,
3'h7,
3'h5,
3'h5,
3'h5,
3'h5,
3'h5,
3'h5,
3'h5,
3'h5,
3'h5,
3'h5,
3'h5,
3'h5,
3'h5,
3'h5,
3'h5,
3'h5,
3'h5,
3'h5,
3'h5,
3'h5,
3'h5,
3'h5,
3'h5,
3'h5,
3'h5,
3'h5,
3'h5,
3'h5,
3'h5,
3'h5,
3'h5,
3'h5,
3'h5,
3'h5,
3'h5,
3'h5,
3'h5,
3'h5,
3'h5,
3'h5,
3'h5,
3'h5,
3'h5,
3'h5,
3'h5,
3'h5,
3'h5,
3'h5,
3'h5,
3'h5,
3'h5,
3'h7,
3'h7,
3'h5,
3'h5,
3'h5,
3'h5,
3'h7,
3'h7,
3'h7,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h7,
3'h0,
3'h0,
3'h0,
3'h7,
3'h7,
3'h0,
3'h0,
3'h7,
3'h0,
3'h7,
3'h7,
3'h0,
3'h7,
3'h7,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h6,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h6,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h6,
3'h0,
3'h0,
3'h0,
3'h6,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h6,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h6,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h6,
3'h6,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h6,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h6,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h6,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h6,
3'h0,
3'h0,
3'h0,
3'h6,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h6,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h6,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h6,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h6,
3'h0,
3'h0,
3'h0,
3'h0,
3'h6,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h6,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h6,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h6,
3'h0,
3'h0,
3'h0,
3'h6,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h6,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h6,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h6,
3'h0,
3'h0,
3'h0,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h0,
3'h0,
3'h6,
3'h6,
3'h6,
3'h6,
3'h0,
3'h0,
3'h6,
3'h6,
3'h0,
3'h0,
3'h6,
3'h0,
3'h0,
3'h6,
3'h6,
3'h6,
3'h0,
3'h0,
3'h6,
3'h0,
3'h6,
3'h6,
3'h6,
3'h0,
3'h6,
3'h6,
3'h6,
3'h0,
3'h0,
3'h6,
3'h6,
3'h0,
3'h0,
3'h6,
3'h0,
3'h6,
3'h6,
3'h0,
3'h0,
3'h6,
3'h6,
3'h0,
3'h6,
3'h6,
3'h0,
3'h0,
3'h6,
3'h6,
3'h0,
3'h0,
3'h6,
3'h0,
3'h0,
3'h6,
3'h6,
3'h0,
3'h6,
3'h6,
3'h0,
3'h6,
3'h0,
3'h0,
3'h0,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h0,
3'h6,
3'h6,
3'h6,
3'h6,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h6,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h6,
3'h6,
3'h6,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h6,
3'h6,
3'h6,
3'h0,
3'h0,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h0,
3'h6,
3'h6,
3'h6,
3'h0,
3'h0,
3'h6,
3'h6,
3'h0,
3'h0,
3'h6,
3'h6,
3'h6,
3'h0,
3'h0,
3'h0,
3'h6,
3'h0,
3'h0,
3'h0,
3'h0,
3'h6,
3'h6,
3'h6,
3'h0,
3'h6,
3'h6,
3'h6,
3'h6,
3'h0,
3'h0,
3'h6,
3'h6,
3'h6,
3'h0,
3'h6,
3'h6,
3'h0,
3'h0,
3'h0,
3'h6,
3'h6,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h6,
3'h0,
3'h0,
3'h6,
3'h0,
3'h7,
3'h0,
3'h7,
3'h0,
3'h0,
3'h0,
3'h7,
3'h7,
3'h7,
3'h0,
3'h0,
3'h7,
3'h7,
3'h7,
3'h7,
3'h0,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h0,
3'h7,
3'h7,
3'h7,
3'h5,
3'h5,
3'h7,
3'h5,
3'h5,
3'h5,
3'h7,
3'h5,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h5,
3'h5,
3'h5,
3'h5,
3'h5,
3'h5,
3'h5,
3'h5,
3'h7,
3'h7,
3'h7,
3'h5,
3'h5,
3'h7,
3'h7,
3'h5,
3'h5,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h5,
3'h7,
3'h7,
3'h5,
3'h5,
3'h7,
3'h7,
3'h5,
3'h7,
3'h5,
3'h5,
3'h7,
3'h7,
3'h5,
3'h5,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h5,
3'h5,
3'h7,
3'h5,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h7,
3'h7,
3'h0,
3'h7,
3'h7,
3'h7,
3'h5,
3'h0,
3'h7,
3'h7,
3'h7,
3'h0,
3'h0,
3'h7,
3'h7,
3'h0,
3'h0,
3'h0,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h0,
3'h7,
3'h7,
3'h0,
3'h0,
3'h6,
3'h0,
3'h0,
3'h6,
3'h6,
3'h0,
3'h0,
3'h0,
3'h0,
3'h6,
3'h6,
3'h0,
3'h0,
3'h0,
3'h6,
3'h0,
3'h6,
3'h6,
3'h0,
3'h0,
3'h6,
3'h6,
3'h6,
3'h0,
3'h0,
3'h0,
3'h6,
3'h6,
3'h0,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h0,
3'h0,
3'h6,
3'h6,
3'h6,
3'h6,
3'h0,
3'h0,
3'h6,
3'h6,
3'h0,
3'h0,
3'h6,
3'h0,
3'h0,
3'h6,
3'h6,
3'h6,
3'h0,
3'h0,
3'h6,
3'h0,
3'h6,
3'h6,
3'h6,
3'h0,
3'h6,
3'h6,
3'h6,
3'h0,
3'h0,
3'h6,
3'h6,
3'h0,
3'h0,
3'h6,
3'h0,
3'h6,
3'h6,
3'h0,
3'h0,
3'h6,
3'h6,
3'h0,
3'h6,
3'h6,
3'h0,
3'h0,
3'h6,
3'h6,
3'h0,
3'h0,
3'h6,
3'h0,
3'h0,
3'h6,
3'h6,
3'h0,
3'h6,
3'h6,
3'h6,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h6,
3'h6,
3'h6,
3'h0,
3'h6,
3'h6,
3'h0,
3'h0,
3'h6,
3'h6,
3'h0,
3'h6,
3'h0,
3'h0,
3'h6,
3'h6,
3'h6,
3'h0,
3'h6,
3'h0,
3'h0,
3'h6,
3'h6,
3'h0,
3'h0,
3'h6,
3'h0,
3'h0,
3'h6,
3'h0,
3'h6,
3'h6,
3'h6,
3'h6,
3'h0,
3'h0,
3'h0,
3'h6,
3'h6,
3'h0,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h0,
3'h0,
3'h6,
3'h6,
3'h6,
3'h6,
3'h0,
3'h0,
3'h6,
3'h6,
3'h0,
3'h0,
3'h6,
3'h0,
3'h0,
3'h6,
3'h6,
3'h6,
3'h0,
3'h0,
3'h6,
3'h0,
3'h6,
3'h6,
3'h6,
3'h0,
3'h6,
3'h6,
3'h6,
3'h0,
3'h0,
3'h6,
3'h6,
3'h0,
3'h0,
3'h6,
3'h0,
3'h6,
3'h6,
3'h0,
3'h0,
3'h6,
3'h6,
3'h0,
3'h6,
3'h6,
3'h0,
3'h0,
3'h6,
3'h6,
3'h0,
3'h0,
3'h6,
3'h0,
3'h0,
3'h6,
3'h6,
3'h0,
3'h6,
3'h6,
3'h0,
3'h6,
3'h6,
3'h6,
3'h6,
3'h0,
3'h6,
3'h6,
3'h0,
3'h6,
3'h6,
3'h6,
3'h0,
3'h6,
3'h6,
3'h0,
3'h6,
3'h6,
3'h0,
3'h0,
3'h6,
3'h6,
3'h0,
3'h6,
3'h0,
3'h6,
3'h6,
3'h0,
3'h6,
3'h6,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h6,
3'h0,
3'h6,
3'h6,
3'h6,
3'h6,
3'h0,
3'h0,
3'h0,
3'h6,
3'h6,
3'h0,
3'h0,
3'h0,
3'h6,
3'h6,
3'h0,
3'h0,
3'h6,
3'h6,
3'h6,
3'h0,
3'h0,
3'h6,
3'h6,
3'h6,
3'h0,
3'h0,
3'h6,
3'h6,
3'h6,
3'h0,
3'h0,
3'h6,
3'h6,
3'h0,
3'h0,
3'h6,
3'h6,
3'h0,
3'h0,
3'h6,
3'h0,
3'h0,
3'h6,
3'h6,
3'h6,
3'h0,
3'h0,
3'h6,
3'h0,
3'h6,
3'h6,
3'h6,
3'h0,
3'h6,
3'h6,
3'h6,
3'h0,
3'h0,
3'h6,
3'h6,
3'h0,
3'h0,
3'h6,
3'h0,
3'h6,
3'h6,
3'h0,
3'h0,
3'h6,
3'h6,
3'h0,
3'h6,
3'h6,
3'h0,
3'h0,
3'h6,
3'h6,
3'h0,
3'h0,
3'h6,
3'h0,
3'h0,
3'h6,
3'h6,
3'h0,
3'h6,
3'h6,
3'h0,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h0,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h6,
3'h6,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h0,
3'h0,
3'h0,
3'h7,
3'h7,
3'h7,
3'h7,
3'h0,
3'h0,
3'h7,
3'h7,
3'h7,
3'h0,
3'h5,
3'h5,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h5,
3'h5,
3'h5,
3'h5,
3'h7,
3'h7,
3'h7,
3'h5,
3'h5,
3'h5,
3'h5,
3'h5,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h5,
3'h5,
3'h5,
3'h7,
3'h7,
3'h7,
3'h5,
3'h5,
3'h5,
3'h7,
3'h7,
3'h7,
3'h7,
3'h0,
3'h0,
3'h0,
3'h7,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h7,
3'h7,
3'h0,
3'h0,
3'h0,
3'h7,
3'h0,
3'h7,
3'h7,
3'h7,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h6,
3'h6,
3'h6,
3'h0,
3'h0,
3'h0,
3'h0,
3'h6,
3'h0,
3'h0,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h0,
3'h6,
3'h6,
3'h6,
3'h6,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h7,
3'h7,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h7,
3'h7,
3'h7,
3'h5,
3'h5,
3'h7,
3'h7,
3'h5,
3'h5,
3'h5,
3'h5,
3'h5,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h5,
3'h5,
3'h5,
3'h5,
3'h7,
3'h7,
3'h5,
3'h5,
3'h5,
3'h7,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h7,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h6,
3'h6,
3'h6,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h6,
3'h0,
3'h6,
3'h0,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h6,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h6,
3'h0,
3'h0,
3'h6,
3'h6,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h6,
3'h6,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h7,
3'h7,
3'h0,
3'h0,
3'h7,
3'h7,
3'h5,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h5,
3'h5,
3'h5,
3'h5,
3'h5,
3'h5,
3'h5,
3'h5,
3'h5,
3'h5,
3'h5,
3'h5,
3'h5,
3'h5,
3'h5,
3'h5,
3'h5,
3'h5,
3'h5,
3'h5,
3'h5,
3'h5,
3'h5,
3'h5,
3'h5,
3'h5,
3'h5,
3'h5,
3'h5,
3'h5,
3'h5,
3'h5,
3'h5,
3'h5,
3'h5,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h0,
3'h0,
3'h0,
3'h7,
3'h0,
3'h0,
3'h7,
3'h7,
3'h0,
3'h0,
3'h6,
3'h6,
3'h6,
3'h6,
3'h0,
3'h6,
3'h6,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h6,
3'h6,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h0,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h6,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h7,
3'h0,
3'h0,
3'h7,
3'h7,
3'h0,
3'h0,
3'h5,
3'h7,
3'h7,
3'h7,
3'h5,
3'h5,
3'h5,
3'h5,
3'h5,
3'h5,
3'h5,
3'h5,
3'h5,
3'h5,
3'h5,
3'h5,
3'h5,
3'h5,
3'h5,
3'h5,
3'h5,
3'h5,
3'h5,
3'h5,
3'h5,
3'h5,
3'h5,
3'h5,
3'h5,
3'h5,
3'h5,
3'h5,
3'h5,
3'h5,
3'h5,
3'h5,
3'h5,
3'h5,
3'h5,
3'h5,
3'h5,
3'h5,
3'h5,
3'h7,
3'h7,
3'h7,
3'h7,
3'h0,
3'h0,
3'h7,
3'h7,
3'h7,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h0,
3'h7,
3'h7,
3'h7,
3'h0,
3'h0,
3'h7,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h5,
3'h0,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h5,
3'h5,
3'h5,
3'h5,
3'h5,
3'h5,
3'h5,
3'h5,
3'h5,
3'h5,
3'h5,
3'h5,
3'h5,
3'h5,
3'h5,
3'h5,
3'h5,
3'h5,
3'h5,
3'h5,
3'h5,
3'h5,
3'h5,
3'h5,
3'h5,
3'h5,
3'h5,
3'h5,
3'h5,
3'h5,
3'h5,
3'h5,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h7,
3'h7,
3'h5,
3'h5,
3'h5,
3'h0,
3'h5,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h6,
3'h6,
3'h0,
3'h0,
3'h0,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h6,
3'h6,
3'h0,
3'h6,
3'h6,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h7,
3'h0,
3'h0,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h0,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h5,
3'h5,
3'h5,
3'h5,
3'h5,
3'h5,
3'h5,
3'h5,
3'h5,
3'h5,
3'h5,
3'h5,
3'h5,
3'h5,
3'h5,
3'h5,
3'h5,
3'h5,
3'h5,
3'h5,
3'h5,
3'h5,
3'h5,
3'h5,
3'h5,
3'h5,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h0,
3'h0,
3'h7,
3'h7,
3'h0,
3'h0,
3'h0,
3'h0,
3'h7,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h6,
3'h6,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h0,
3'h6,
3'h6,
3'h6,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h6,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h6,
3'h6,
3'h0,
3'h0,
3'h0,
3'h7,
3'h7,
3'h0,
3'h7,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h7,
3'h5,
3'h5,
3'h0,
3'h0,
3'h5,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h5,
3'h5,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h6,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h6,
3'h6,
3'h0,
3'h0,
3'h6,
3'h0,
3'h0,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h0,
3'h0,
3'h6,
3'h6,
3'h6,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h7,
3'h0,
3'h0,
3'h7,
3'h7,
3'h0,
3'h7,
3'h7,
3'h0,
3'h0,
3'h7,
3'h7,
3'h7,
3'h0,
3'h0,
3'h0,
3'h0,
3'h5,
3'h7,
3'h7,
3'h5,
3'h5,
3'h5,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h5,
3'h5,
3'h5,
3'h5,
3'h5,
3'h5,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h7,
3'h0,
3'h0,
3'h0,
3'h7,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h7,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h6,
3'h0,
3'h0,
3'h0,
3'h6,
3'h0,
3'h0,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h7,
3'h7,
3'h7,
3'h5,
3'h0,
3'h7,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h7,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h7,
3'h7,
3'h7,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h7,
3'h0,
3'h0,
3'h0,
3'h0,
3'h7,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h6,
3'h0,
3'h0,
3'h0,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h6,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h6,
3'h6,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h6,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h0,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h0,
3'h0,
3'h0,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h0,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h0,
3'h6,
3'h6,
3'h0,
3'h0,
3'h6,
3'h6,
3'h6,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h6,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h6,
3'h0,
3'h0,
3'h0,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h0,
3'h0,
3'h6,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h0,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h0,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h0,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h0,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h0,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h0,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h1,
3'h1,
3'h1,
3'h1,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h1,
3'h1,
3'h1,
3'h1,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h1,
3'h1,
3'h1,
3'h1,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h1,
3'h1,
3'h6,
3'h1,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h1,
3'h1,
3'h6,
3'h1,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h1,
3'h1,
3'h1,
3'h1,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h1,
3'h1,
3'h1,
3'h1,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h1,
3'h1,
3'h4,
3'h1,
3'h5,
3'h1,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h1,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h1,
3'h1,
3'h4,
3'h1,
3'h5,
3'h1,
3'h1,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h1,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h1,
3'h1,
3'h5,
3'h1,
3'h4,
3'h1,
3'h1,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h1,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h1,
3'h5,
3'h1,
3'h1,
3'h5,
3'h1,
3'h1,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h0,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h1,
3'h5,
3'h1,
3'h1,
3'h5,
3'h1,
3'h1,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h0,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h1,
3'h1,
3'h4,
3'h1,
3'h5,
3'h1,
3'h1,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h1,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h1,
3'h1,
3'h5,
3'h1,
3'h4,
3'h1,
3'h1,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h1,
3'h1,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h1,
3'h1,
3'h1,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h1,
3'h1,
3'h5,
3'h1,
3'h4,
3'h4,
3'h1,
3'h4,
3'h1,
3'h1,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h1,
3'h1,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h1,
3'h1,
3'h1,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h1,
3'h5,
3'h1,
3'h4,
3'h4,
3'h1,
3'h4,
3'h1,
3'h1,
3'h1,
3'h1,
3'h6,
3'h1,
3'h6,
3'h1,
3'h6,
3'h1,
3'h1,
3'h1,
3'h6,
3'h6,
3'h6,
3'h1,
3'h1,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h1,
3'h1,
3'h1,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h1,
3'h1,
3'h1,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h1,
3'h6,
3'h1,
3'h1,
3'h4,
3'h1,
3'h4,
3'h4,
3'h1,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h6,
3'h6,
3'h6,
3'h1,
3'h1,
3'h0,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h1,
3'h1,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h1,
3'h1,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h1,
3'h1,
3'h1,
3'h1,
3'h4,
3'h1,
3'h1,
3'h5,
3'h1,
3'h1,
3'h1,
3'h1,
3'h6,
3'h6,
3'h6,
3'h1,
3'h1,
3'h1,
3'h1,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h1,
3'h1,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h1,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h1,
3'h1,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h1,
3'h1,
3'h1,
3'h1,
3'h4,
3'h1,
3'h1,
3'h5,
3'h1,
3'h1,
3'h1,
3'h1,
3'h6,
3'h6,
3'h6,
3'h1,
3'h1,
3'h1,
3'h1,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h1,
3'h1,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h1,
3'h1,
3'h1,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h1,
3'h5,
3'h1,
3'h4,
3'h4,
3'h1,
3'h4,
3'h1,
3'h1,
3'h1,
3'h1,
3'h6,
3'h1,
3'h6,
3'h1,
3'h6,
3'h6,
3'h1,
3'h1,
3'h6,
3'h6,
3'h1,
3'h1,
3'h1,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h1,
3'h1,
3'h1,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h1,
3'h1,
3'h1,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h1,
3'h6,
3'h1,
3'h1,
3'h4,
3'h1,
3'h4,
3'h4,
3'h1,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h1,
3'h1,
3'h6,
3'h1,
3'h1,
3'h6,
3'h6,
3'h6,
3'h1,
3'h1,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h1,
3'h1,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h1,
3'h1,
3'h5,
3'h1,
3'h1,
3'h6,
3'h6,
3'h1,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h1,
3'h6,
3'h1,
3'h1,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h1,
3'h5,
3'h5,
3'h1,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h0,
3'h1,
3'h1,
3'h4,
3'h1,
3'h1,
3'h6,
3'h1,
3'h6,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h5,
3'h1,
3'h4,
3'h4,
3'h4,
3'h1,
3'h4,
3'h4,
3'h5,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h6,
3'h1,
3'h1,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h1,
3'h5,
3'h5,
3'h1,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h0,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h0,
3'h1,
3'h1,
3'h4,
3'h1,
3'h6,
3'h6,
3'h6,
3'h6,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h5,
3'h1,
3'h4,
3'h4,
3'h1,
3'h1,
3'h4,
3'h4,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h5,
3'h1,
3'h1,
3'h5,
3'h1,
3'h1,
3'h1,
3'h1,
3'h5,
3'h1,
3'h1,
3'h6,
3'h6,
3'h1,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h1,
3'h6,
3'h6,
3'h1,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h1,
3'h1,
3'h4,
3'h1,
3'h6,
3'h6,
3'h1,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h1,
3'h1,
3'h5,
3'h1,
3'h1,
3'h6,
3'h6,
3'h6,
3'h6,
3'h1,
3'h1,
3'h1,
3'h1,
3'h5,
3'h1,
3'h1,
3'h4,
3'h4,
3'h1,
3'h4,
3'h4,
3'h5,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h5,
3'h5,
3'h1,
3'h5,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h5,
3'h1,
3'h6,
3'h6,
3'h6,
3'h1,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h1,
3'h6,
3'h1,
3'h6,
3'h6,
3'h6,
3'h1,
3'h6,
3'h6,
3'h1,
3'h5,
3'h1,
3'h1,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h1,
3'h4,
3'h4,
3'h1,
3'h6,
3'h6,
3'h6,
3'h6,
3'h1,
3'h1,
3'h1,
3'h1,
3'h5,
3'h1,
3'h1,
3'h5,
3'h4,
3'h1,
3'h4,
3'h4,
3'h4,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h5,
3'h1,
3'h5,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h5,
3'h1,
3'h1,
3'h6,
3'h6,
3'h1,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h1,
3'h6,
3'h1,
3'h1,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h1,
3'h5,
3'h5,
3'h1,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h1,
3'h1,
3'h5,
3'h1,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h1,
3'h4,
3'h4,
3'h1,
3'h6,
3'h6,
3'h6,
3'h6,
3'h1,
3'h1,
3'h1,
3'h1,
3'h5,
3'h1,
3'h1,
3'h5,
3'h4,
3'h1,
3'h4,
3'h4,
3'h4,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h5,
3'h1,
3'h5,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h5,
3'h1,
3'h1,
3'h6,
3'h6,
3'h1,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h1,
3'h6,
3'h1,
3'h1,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h1,
3'h5,
3'h5,
3'h1,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h0,
3'h1,
3'h1,
3'h4,
3'h1,
3'h1,
3'h6,
3'h1,
3'h6,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h5,
3'h1,
3'h4,
3'h4,
3'h1,
3'h1,
3'h4,
3'h4,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h5,
3'h1,
3'h1,
3'h5,
3'h1,
3'h1,
3'h1,
3'h1,
3'h5,
3'h1,
3'h1,
3'h6,
3'h6,
3'h1,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h1,
3'h6,
3'h6,
3'h1,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h1,
3'h1,
3'h5,
3'h1,
3'h6,
3'h6,
3'h1,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h1,
3'h1,
3'h4,
3'h1,
3'h1,
3'h6,
3'h1,
3'h6,
3'h6,
3'h1,
3'h1,
3'h1,
3'h1,
3'h5,
3'h1,
3'h1,
3'h4,
3'h4,
3'h1,
3'h4,
3'h4,
3'h5,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h5,
3'h5,
3'h1,
3'h5,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h5,
3'h1,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h1,
3'h6,
3'h6,
3'h6,
3'h1,
3'h6,
3'h6,
3'h1,
3'h5,
3'h1,
3'h1,
3'h6,
3'h1,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h1,
3'h1,
3'h4,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h6,
3'h6,
3'h6,
3'h6,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h6,
3'h6,
3'h1,
3'h1,
3'h1,
3'h1,
3'h4,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h1,
3'h1,
3'h4,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h4,
3'h4,
3'h1,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h6,
3'h6,
3'h1,
3'h1,
3'h1,
3'h1,
3'h4,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h1,
3'h1,
3'h4,
3'h1,
3'h1,
3'h6,
3'h6,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h4,
3'h4,
3'h1,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h5,
3'h4,
3'h1,
3'h4,
3'h1,
3'h1,
3'h1,
3'h1,
3'h4,
3'h1,
3'h1,
3'h1,
3'h6,
3'h1,
3'h1,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h6,
3'h6,
3'h6,
3'h1,
3'h1,
3'h1,
3'h4,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h1,
3'h1,
3'h4,
3'h1,
3'h1,
3'h1,
3'h1,
3'h6,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h4,
3'h1,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h4,
3'h4,
3'h1,
3'h4,
3'h1,
3'h1,
3'h1,
3'h1,
3'h4,
3'h1,
3'h1,
3'h6,
3'h6,
3'h6,
3'h1,
3'h1,
3'h6,
3'h6,
3'h6,
3'h6,
3'h1,
3'h1,
3'h1,
3'h1,
3'h6,
3'h6,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h4,
3'h1,
3'h1,
3'h1,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h1,
3'h1,
3'h1,
3'h4,
3'h4,
3'h1,
3'h1,
3'h6,
3'h6,
3'h6,
3'h1,
3'h1,
3'h1,
3'h1,
3'h4,
3'h1,
3'h1,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h5,
3'h1,
3'h4,
3'h4,
3'h1,
3'h1,
3'h1,
3'h1,
3'h4,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h6,
3'h6,
3'h6,
3'h6,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h6,
3'h6,
3'h1,
3'h1,
3'h1,
3'h1,
3'h4,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h0,
3'h1,
3'h1,
3'h1,
3'h4,
3'h1,
3'h1,
3'h0,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h1,
3'h1,
3'h1,
3'h4,
3'h4,
3'h1,
3'h1,
3'h6,
3'h6,
3'h6,
3'h1,
3'h1,
3'h1,
3'h1,
3'h4,
3'h1,
3'h1,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h5,
3'h1,
3'h4,
3'h4,
3'h1,
3'h1,
3'h1,
3'h1,
3'h4,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h6,
3'h6,
3'h6,
3'h6,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h6,
3'h6,
3'h1,
3'h1,
3'h1,
3'h1,
3'h4,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h1,
3'h1,
3'h4,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h4,
3'h4,
3'h1,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h5,
3'h1,
3'h1,
3'h4,
3'h1,
3'h1,
3'h1,
3'h1,
3'h4,
3'h1,
3'h1,
3'h6,
3'h6,
3'h1,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h6,
3'h6,
3'h6,
3'h1,
3'h1,
3'h1,
3'h4,
3'h1,
3'h1,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h1,
3'h1,
3'h4,
3'h1,
3'h1,
3'h1,
3'h1,
3'h6,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h4,
3'h1,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h5,
3'h4,
3'h1,
3'h4,
3'h1,
3'h1,
3'h1,
3'h1,
3'h4,
3'h1,
3'h1,
3'h1,
3'h6,
3'h6,
3'h1,
3'h1,
3'h6,
3'h6,
3'h6,
3'h6,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h4,
3'h1,
3'h1,
3'h1,
3'h1,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h4,
3'h4,
3'h4,
3'h4,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h5,
3'h1,
3'h4,
3'h4,
3'h1,
3'h1,
3'h4,
3'h4,
3'h1,
3'h5,
3'h4,
3'h4,
3'h5,
3'h1,
3'h4,
3'h1,
3'h1,
3'h6,
3'h6,
3'h6,
3'h6,
3'h1,
3'h6,
3'h6,
3'h1,
3'h6,
3'h1,
3'h1,
3'h1,
3'h1,
3'h6,
3'h6,
3'h1,
3'h0,
3'h6,
3'h1,
3'h1,
3'h1,
3'h4,
3'h4,
3'h4,
3'h4,
3'h1,
3'h1,
3'h5,
3'h1,
3'h1,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h5,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h4,
3'h1,
3'h1,
3'h5,
3'h4,
3'h4,
3'h5,
3'h1,
3'h4,
3'h1,
3'h1,
3'h6,
3'h6,
3'h6,
3'h6,
3'h1,
3'h6,
3'h6,
3'h1,
3'h6,
3'h1,
3'h1,
3'h1,
3'h1,
3'h6,
3'h6,
3'h1,
3'h0,
3'h6,
3'h1,
3'h1,
3'h1,
3'h4,
3'h4,
3'h4,
3'h4,
3'h1,
3'h1,
3'h5,
3'h1,
3'h1,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h1,
3'h1,
3'h5,
3'h5,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h5,
3'h1,
3'h1,
3'h5,
3'h1,
3'h1,
3'h1,
3'h5,
3'h1,
3'h4,
3'h4,
3'h4,
3'h4,
3'h1,
3'h1,
3'h4,
3'h1,
3'h1,
3'h6,
3'h6,
3'h6,
3'h1,
3'h1,
3'h0,
3'h1,
3'h6,
3'h6,
3'h1,
3'h1,
3'h1,
3'h1,
3'h0,
3'h1,
3'h6,
3'h6,
3'h1,
3'h1,
3'h1,
3'h1,
3'h4,
3'h4,
3'h4,
3'h4,
3'h1,
3'h5,
3'h1,
3'h1,
3'h5,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h5,
3'h1,
3'h1,
3'h1,
3'h5,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h4,
3'h1,
3'h5,
3'h1,
3'h1,
3'h1,
3'h5,
3'h1,
3'h1,
3'h4,
3'h4,
3'h4,
3'h1,
3'h1,
3'h5,
3'h1,
3'h1,
3'h0,
3'h6,
3'h6,
3'h6,
3'h1,
3'h6,
3'h6,
3'h1,
3'h6,
3'h1,
3'h1,
3'h1,
3'h1,
3'h6,
3'h6,
3'h6,
3'h6,
3'h1,
3'h1,
3'h1,
3'h1,
3'h4,
3'h4,
3'h4,
3'h4,
3'h1,
3'h5,
3'h1,
3'h1,
3'h5,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h5,
3'h1,
3'h4,
3'h4,
3'h1,
3'h1,
3'h4,
3'h4,
3'h1,
3'h5,
3'h4,
3'h4,
3'h5,
3'h1,
3'h4,
3'h1,
3'h1,
3'h6,
3'h6,
3'h6,
3'h6,
3'h1,
3'h6,
3'h6,
3'h1,
3'h6,
3'h1,
3'h1,
3'h1,
3'h1,
3'h6,
3'h6,
3'h1,
3'h0,
3'h6,
3'h1,
3'h1,
3'h1,
3'h4,
3'h4,
3'h4,
3'h4,
3'h1,
3'h1,
3'h0,
3'h6,
3'h6,
3'h6,
3'h1,
3'h6,
3'h6,
3'h1,
3'h6,
3'h1,
3'h1,
3'h1,
3'h1,
3'h6,
3'h6,
3'h6,
3'h6,
3'h1,
3'h1,
3'h1,
3'h1,
3'h4,
3'h4,
3'h4,
3'h4,
3'h1,
3'h5,
3'h1,
3'h1,
3'h5,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h5,
3'h1,
3'h4,
3'h4,
3'h1,
3'h1,
3'h4,
3'h4,
3'h1,
3'h5,
3'h4,
3'h4,
3'h5,
3'h1,
3'h4,
3'h1,
3'h1,
3'h6,
3'h6,
3'h6,
3'h6,
3'h1,
3'h6,
3'h6,
3'h1,
3'h6,
3'h1,
3'h1,
3'h1,
3'h1,
3'h6,
3'h6,
3'h1,
3'h0,
3'h6,
3'h1,
3'h1,
3'h1,
3'h4,
3'h4,
3'h4,
3'h4,
3'h1,
3'h1,
3'h5,
3'h1,
3'h1,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h1,
3'h1,
3'h5,
3'h5,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h5,
3'h1,
3'h1,
3'h5,
3'h1,
3'h1,
3'h1,
3'h5,
3'h1,
3'h1,
3'h4,
3'h4,
3'h4,
3'h1,
3'h1,
3'h5,
3'h1,
3'h1,
3'h6,
3'h6,
3'h6,
3'h6,
3'h6,
3'h0,
3'h1,
3'h6,
3'h6,
3'h1,
3'h1,
3'h1,
3'h1,
3'h0,
3'h1,
3'h6,
3'h6,
3'h1,
3'h1,
3'h1,
3'h1,
3'h4,
3'h4,
3'h4,
3'h1,
3'h1,
3'h5,
3'h1,
3'h1,
3'h5,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h5,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h5,
3'h1,
3'h1,
3'h1,
3'h3,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h5,
3'h1,
3'h5,
3'h1,
3'h1,
3'h1,
3'h5,
3'h1,
3'h1,
3'h4,
3'h4,
3'h4,
3'h1,
3'h1,
3'h5,
3'h1,
3'h1,
3'h0,
3'h6,
3'h6,
3'h6,
3'h1,
3'h6,
3'h4,
3'h4,
3'h4,
3'h4,
3'h1,
3'h1,
3'h1,
3'h5,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h4,
3'h4,
3'h1,
3'h4,
3'h4,
3'h1,
3'h4,
3'h4,
3'h4,
3'h1,
3'h4,
3'h4,
3'h4,
3'h4,
3'h1,
3'h4,
3'h4,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h1,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h1,
3'h4,
3'h4,
3'h1,
3'h1,
3'h4,
3'h4,
3'h1,
3'h4,
3'h4,
3'h4,
3'h4,
3'h1,
3'h4,
3'h4,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h4,
3'h1,
3'h4,
3'h4,
3'h4,
3'h4,
3'h1,
3'h4,
3'h4,
3'h1,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h1,
3'h4,
3'h1,
3'h4,
3'h4,
3'h1,
3'h4,
3'h1,
3'h4,
3'h1,
3'h4,
3'h1,
3'h4,
3'h4,
3'h1,
3'h1,
3'h1,
3'h4,
3'h1,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h1,
3'h4,
3'h1,
3'h1,
3'h1,
3'h6,
3'h6,
3'h6,
3'h1,
3'h1,
3'h1,
3'h6,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h5,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h1,
3'h1,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h1,
3'h1,
3'h1,
3'h4,
3'h4,
3'h1,
3'h1,
3'h1,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h1,
3'h4,
3'h1,
3'h4,
3'h1,
3'h1,
3'h4,
3'h4,
3'h4,
3'h4,
3'h1,
3'h4,
3'h4,
3'h1,
3'h1,
3'h6,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h4,
3'h4,
3'h4,
3'h4,
3'h1,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h1,
3'h1,
3'h1,
3'h5,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h4,
3'h4,
3'h1,
3'h4,
3'h4,
3'h1,
3'h4,
3'h4,
3'h4,
3'h1,
3'h4,
3'h4,
3'h4,
3'h4,
3'h1,
3'h4,
3'h4,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h4,
3'h1,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h1,
3'h1,
3'h6,
3'h1,
3'h1,
3'h0,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h4,
3'h4,
3'h4,
3'h4,
3'h1,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h1,
3'h1,
3'h1,
3'h5,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h4,
3'h4,
3'h1,
3'h4,
3'h4,
3'h1,
3'h4,
3'h4,
3'h4,
3'h1,
3'h4,
3'h4,
3'h4,
3'h4,
3'h1,
3'h4,
3'h4,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h1,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h1,
3'h1,
3'h1,
3'h4,
3'h1,
3'h4,
3'h1,
3'h4,
3'h4,
3'h1,
3'h1,
3'h4,
3'h4,
3'h1,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h1,
3'h4,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h1,
3'h4,
3'h4,
3'h4,
3'h1,
3'h1,
3'h1,
3'h1,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h1,
3'h4,
3'h1,
3'h4,
3'h4,
3'h1,
3'h4,
3'h4,
3'h4,
3'h4,
3'h1,
3'h4,
3'h4,
3'h1,
3'h1,
3'h6,
3'h1,
3'h1,
3'h1,
3'h1,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h5,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h1,
3'h1,
3'h1,
3'h1,
3'h5,
3'h1,
3'h1,
3'h5,
3'h1,
3'h1,
3'h4,
3'h4,
3'h5,
3'h1,
3'h1,
3'h5,
3'h1,
3'h1,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h1,
3'h1,
3'h1,
3'h1,
3'h5,
3'h1,
3'h1,
3'h4,
3'h1,
3'h1,
3'h4,
3'h4,
3'h4,
3'h1,
3'h1,
3'h3,
3'h1,
3'h1,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h1,
3'h1,
3'h1,
3'h1,
3'h5,
3'h4,
3'h1,
3'h3,
3'h1,
3'h1,
3'h4,
3'h4,
3'h4,
3'h4,
3'h1,
3'h5,
3'h1,
3'h1,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h1,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h1,
3'h1,
3'h1,
3'h1,
3'h5,
3'h1,
3'h1,
3'h4,
3'h1,
3'h4,
3'h4,
3'h4,
3'h4,
3'h1,
3'h4,
3'h4,
3'h1,
3'h5,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h5,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h1,
3'h1,
3'h1,
3'h1,
3'h5,
3'h1,
3'h1,
3'h5,
3'h1,
3'h1,
3'h4,
3'h4,
3'h5,
3'h1,
3'h1,
3'h5,
3'h1,
3'h1,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h1,
3'h1,
3'h1,
3'h1,
3'h5,
3'h1,
3'h1,
3'h4,
3'h1,
3'h4,
3'h4,
3'h4,
3'h4,
3'h1,
3'h4,
3'h4,
3'h1,
3'h5,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h5,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h1,
3'h1,
3'h1,
3'h1,
3'h5,
3'h1,
3'h1,
3'h5,
3'h1,
3'h1,
3'h4,
3'h4,
3'h5,
3'h1,
3'h1,
3'h5,
3'h1,
3'h1,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h1,
3'h1,
3'h1,
3'h1,
3'h5,
3'h1,
3'h1,
3'h5,
3'h1,
3'h1,
3'h4,
3'h4,
3'h4,
3'h1,
3'h1,
3'h5,
3'h1,
3'h1,
3'h5,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h1,
3'h1,
3'h1,
3'h1,
3'h5,
3'h1,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h1,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h1,
3'h5,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h1,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h1,
3'h4,
3'h4,
3'h4,
3'h1,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h1,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h1,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h1,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h1,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h1,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h1,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h1,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h1,
3'h4,
3'h4,
3'h1,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h1,
3'h1,
3'h4,
3'h1,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h1,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h1,
3'h4,
3'h4,
3'h1,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h1,
3'h4,
3'h1,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h1,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h1,
3'h4,
3'h4,
3'h1,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h1,
3'h4,
3'h4,
3'h1,
3'h4,
3'h1,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h1,
3'h1,
3'h4,
3'h1,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h1,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h1,
3'h1,
3'h4,
3'h1,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h1,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h1,
3'h4,
3'h1,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h1,
3'h4,
3'h1,
3'h4,
3'h4,
3'h1,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h1,
3'h4,
3'h4,
3'h1,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h1,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h1,
3'h4,
3'h1,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h1,
3'h4,
3'h4,
3'h1,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h1,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h1,
3'h4,
3'h1,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h1,
3'h4,
3'h1,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h1,
3'h1,
3'h4,
3'h1,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h1,
3'h1,
3'h4,
3'h1,
3'h4,
3'h4,
3'h1,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h1,
3'h1,
3'h4,
3'h1,
3'h4,
3'h4,
3'h1,
3'h4,
3'h4,
3'h1,
3'h4,
3'h1,
3'h4,
3'h4,
3'h1,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h1,
3'h4,
3'h1,
3'h1,
3'h4,
3'h1,
3'h4,
3'h4,
3'h1,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h1,
3'h4,
3'h4,
3'h4,
3'h4,
3'h1,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h1,
3'h4,
3'h1,
3'h1,
3'h4,
3'h1,
3'h4,
3'h4,
3'h1,
3'h4,
3'h4,
3'h4,
3'h1,
3'h4,
3'h1,
3'h1,
3'h4,
3'h1,
3'h4,
3'h4,
3'h1,
3'h4,
3'h4,
3'h4,
3'h4,
3'h1,
3'h4,
3'h4,
3'h1,
3'h4,
3'h1,
3'h1,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h1,
3'h1,
3'h4,
3'h1,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h1,
3'h1,
3'h4,
3'h1,
3'h4,
3'h4,
3'h1,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h1,
3'h1,
3'h4,
3'h1,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h1,
3'h1,
3'h4,
3'h1,
3'h4,
3'h4,
3'h1,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h1,
3'h1,
3'h4,
3'h1,
3'h4,
3'h4,
3'h1,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h1,
3'h1,
3'h4,
3'h1,
3'h4,
3'h4,
3'h1,
3'h4,
3'h4,
3'h4,
3'h4,
3'h1,
3'h4,
3'h4,
3'h1,
3'h4,
3'h1,
3'h1,
3'h4,
3'h1,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h1,
3'h4,
3'h4,
3'h1,
3'h4,
3'h4,
3'h1,
3'h4,
3'h1,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h1,
3'h4,
3'h4,
3'h1,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h1,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h1,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h1,
3'h4,
3'h4,
3'h4,
3'h4,
3'h1,
3'h4,
3'h4,
3'h1,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h1,
3'h4,
3'h4,
3'h1,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h1,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h1,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h1,
3'h4,
3'h4,
3'h4,
3'h4,
3'h1,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h1,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h1,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h1,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h1,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h1,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h1,
3'h4,
3'h4,
3'h1,
3'h4,
3'h4,
3'h1,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h1,
3'h4,
3'h4,
3'h1,
3'h4,
3'h4,
3'h4,
3'h4,
3'h1,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h1,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h1,
3'h4,
3'h4,
3'h1,
3'h4,
3'h4,
3'h1,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h1,
3'h4,
3'h4,
3'h1,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h1,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h1,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h1,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h1,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h1,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h1,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h1,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h1,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h1,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h1,
3'h1,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h1,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h1,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h1,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h1,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h1,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h1,
3'h1,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h1,
3'h1,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h1,
3'h1,
3'h4,
3'h1,
3'h1,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h1,
3'h1,
3'h4,
3'h4,
3'h4,
3'h4,
3'h1,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h1,
3'h1,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h1,
3'h1,
3'h4,
3'h1,
3'h1,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h1,
3'h1,
3'h4,
3'h4,
3'h4,
3'h4,
3'h1,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h1,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h1,
3'h4,
3'h1,
3'h1,
3'h1,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h1,
3'h4,
3'h4,
3'h4,
3'h4,
3'h1,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h1,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h1,
3'h4,
3'h4,
3'h1,
3'h1,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h1,
3'h4,
3'h4,
3'h4,
3'h4,
3'h1,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h1,
3'h1,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h1,
3'h1,
3'h4,
3'h1,
3'h1,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h1,
3'h1,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h1,
3'h4,
3'h4,
3'h1,
3'h1,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h1,
3'h4,
3'h4,
3'h4,
3'h4,
3'h1,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h1,
3'h1,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h1,
3'h1,
3'h4,
3'h1,
3'h1,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h1,
3'h1,
3'h4,
3'h4,
3'h4,
3'h4,
3'h1,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h1,
3'h4,
3'h1,
3'h1,
3'h1,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h1,
3'h4,
3'h4,
3'h4,
3'h4,
3'h1,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h1,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h1,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h1,
3'h1,
3'h4,
3'h1,
3'h4,
3'h4,
3'h4,
3'h1,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h1,
3'h1,
3'h4,
3'h1,
3'h1,
3'h1,
3'h4,
3'h4,
3'h4,
3'h4,
3'h1,
3'h4,
3'h1,
3'h1,
3'h4,
3'h4,
3'h4,
3'h1,
3'h1,
3'h4,
3'h4,
3'h4,
3'h1,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h1,
3'h4,
3'h1,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h1,
3'h1,
3'h4,
3'h1,
3'h1,
3'h1,
3'h4,
3'h4,
3'h4,
3'h4,
3'h1,
3'h4,
3'h1,
3'h1,
3'h4,
3'h4,
3'h4,
3'h1,
3'h1,
3'h4,
3'h4,
3'h4,
3'h1,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h1,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h1,
3'h4,
3'h1,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h1,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h1,
3'h1,
3'h4,
3'h1,
3'h1,
3'h1,
3'h1,
3'h4,
3'h4,
3'h4,
3'h1,
3'h4,
3'h4,
3'h1,
3'h4,
3'h4,
3'h4,
3'h4,
3'h1,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h1,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h1,
3'h1,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h1,
3'h1,
3'h4,
3'h4,
3'h1,
3'h1,
3'h1,
3'h4,
3'h4,
3'h4,
3'h1,
3'h1,
3'h4,
3'h1,
3'h1,
3'h4,
3'h4,
3'h4,
3'h1,
3'h1,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h1,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h1,
3'h1,
3'h4,
3'h1,
3'h4,
3'h4,
3'h4,
3'h1,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h1,
3'h1,
3'h4,
3'h1,
3'h1,
3'h1,
3'h4,
3'h4,
3'h4,
3'h4,
3'h1,
3'h4,
3'h4,
3'h1,
3'h4,
3'h4,
3'h4,
3'h1,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h1,
3'h1,
3'h4,
3'h4,
3'h1,
3'h1,
3'h1,
3'h4,
3'h4,
3'h4,
3'h1,
3'h1,
3'h4,
3'h1,
3'h1,
3'h4,
3'h4,
3'h4,
3'h1,
3'h1,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h1,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h1,
3'h1,
3'h4,
3'h1,
3'h4,
3'h4,
3'h4,
3'h1,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h1,
3'h1,
3'h4,
3'h1,
3'h1,
3'h1,
3'h4,
3'h4,
3'h4,
3'h4,
3'h1,
3'h4,
3'h1,
3'h1,
3'h4,
3'h4,
3'h4,
3'h1,
3'h1,
3'h4,
3'h4,
3'h4,
3'h1,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h1,
3'h1,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h1,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h1,
3'h1,
3'h4,
3'h1,
3'h1,
3'h1,
3'h1,
3'h4,
3'h4,
3'h4,
3'h1,
3'h4,
3'h4,
3'h1,
3'h4,
3'h4,
3'h4,
3'h4,
3'h1,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h1,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h1,
3'h1,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h1,
3'h4,
3'h1,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h1,
3'h4,
3'h4,
3'h4,
3'h1,
3'h1,
3'h1,
3'h4,
3'h1,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h1,
3'h1,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h1,
3'h1,
3'h1,
3'h4,
3'h1,
3'h1,
3'h1,
3'h1,
3'h4,
3'h4,
3'h1,
3'h1,
3'h4,
3'h1,
3'h1,
3'h1,
3'h4,
3'h1,
3'h1,
3'h1,
3'h4,
3'h4,
3'h4,
3'h1,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h1,
3'h4,
3'h4,
3'h4,
3'h1,
3'h4,
3'h4,
3'h4,
3'h1,
3'h1,
3'h1,
3'h4,
3'h1,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h1,
3'h1,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h1,
3'h1,
3'h1,
3'h4,
3'h1,
3'h1,
3'h1,
3'h1,
3'h4,
3'h4,
3'h1,
3'h1,
3'h4,
3'h1,
3'h1,
3'h1,
3'h4,
3'h1,
3'h1,
3'h1,
3'h4,
3'h4,
3'h4,
3'h1,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h1,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h1,
3'h4,
3'h4,
3'h1,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h1,
3'h1,
3'h4,
3'h1,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h1,
3'h1,
3'h1,
3'h4,
3'h1,
3'h1,
3'h1,
3'h1,
3'h4,
3'h4,
3'h4,
3'h1,
3'h1,
3'h4,
3'h1,
3'h1,
3'h4,
3'h4,
3'h1,
3'h1,
3'h1,
3'h4,
3'h4,
3'h1,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h1,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h1,
3'h4,
3'h4,
3'h1,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h1,
3'h4,
3'h4,
3'h4,
3'h1,
3'h1,
3'h4,
3'h4,
3'h1,
3'h4,
3'h4,
3'h4,
3'h1,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h1,
3'h1,
3'h4,
3'h4,
3'h1,
3'h1,
3'h1,
3'h1,
3'h4,
3'h4,
3'h1,
3'h1,
3'h4,
3'h1,
3'h1,
3'h4,
3'h4,
3'h1,
3'h1,
3'h1,
3'h4,
3'h4,
3'h1,
3'h1,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h1,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h1,
3'h4,
3'h1,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h1,
3'h4,
3'h4,
3'h4,
3'h1,
3'h1,
3'h1,
3'h4,
3'h1,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h1,
3'h1,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h1,
3'h1,
3'h1,
3'h4,
3'h1,
3'h1,
3'h1,
3'h1,
3'h4,
3'h4,
3'h4,
3'h1,
3'h4,
3'h1,
3'h1,
3'h1,
3'h4,
3'h4,
3'h4,
3'h1,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h1,
3'h1,
3'h4,
3'h4,
3'h1,
3'h1,
3'h1,
3'h1,
3'h4,
3'h4,
3'h1,
3'h1,
3'h4,
3'h1,
3'h1,
3'h4,
3'h4,
3'h1,
3'h1,
3'h1,
3'h4,
3'h4,
3'h1,
3'h1,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h1,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h1,
3'h4,
3'h1,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h1,
3'h4,
3'h4,
3'h4,
3'h1,
3'h1,
3'h1,
3'h4,
3'h1,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h1,
3'h1,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h1,
3'h1,
3'h1,
3'h4,
3'h1,
3'h1,
3'h1,
3'h1,
3'h4,
3'h4,
3'h1,
3'h1,
3'h4,
3'h1,
3'h1,
3'h1,
3'h4,
3'h1,
3'h1,
3'h1,
3'h4,
3'h4,
3'h4,
3'h1,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h1,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h1,
3'h4,
3'h4,
3'h1,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h1,
3'h4,
3'h4,
3'h4,
3'h1,
3'h1,
3'h4,
3'h1,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h1,
3'h1,
3'h1,
3'h4,
3'h1,
3'h1,
3'h1,
3'h1,
3'h4,
3'h4,
3'h4,
3'h1,
3'h1,
3'h4,
3'h1,
3'h1,
3'h4,
3'h4,
3'h1,
3'h1,
3'h4,
3'h4,
3'h4,
3'h1,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h1,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h1,
3'h4,
3'h4,
3'h1,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h1,
3'h4,
3'h4,
3'h4,
3'h1,
3'h1,
3'h4,
3'h4,
3'h1,
3'h4,
3'h4,
3'h4,
3'h1,
3'h4,
3'h4,
3'h4,
3'h1,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h1,
3'h4,
3'h5,
3'h1,
3'h1,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h1,
3'h4,
3'h4,
3'h4,
3'h1,
3'h4,
3'h4,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h4,
3'h4,
3'h1,
3'h4,
3'h4,
3'h4,
3'h1,
3'h1,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h4,
3'h4,
3'h1,
3'h4,
3'h4,
3'h4,
3'h1,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h1,
3'h1,
3'h4,
3'h4,
3'h1,
3'h4,
3'h4,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h4,
3'h4,
3'h1,
3'h4,
3'h4,
3'h4,
3'h1,
3'h1,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h4,
3'h4,
3'h1,
3'h4,
3'h4,
3'h4,
3'h1,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h1,
3'h1,
3'h4,
3'h4,
3'h1,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h1,
3'h1,
3'h4,
3'h1,
3'h1,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h1,
3'h1,
3'h4,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h4,
3'h4,
3'h1,
3'h1,
3'h4,
3'h4,
3'h1,
3'h1,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h4,
3'h1,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h1,
3'h1,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h1,
3'h4,
3'h4,
3'h1,
3'h1,
3'h4,
3'h4,
3'h1,
3'h4,
3'h4,
3'h4,
3'h1,
3'h4,
3'h4,
3'h4,
3'h1,
3'h4,
3'h4,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h4,
3'h4,
3'h1,
3'h4,
3'h4,
3'h4,
3'h1,
3'h1,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h4,
3'h1,
3'h1,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h1,
3'h4,
3'h4,
3'h1,
3'h1,
3'h4,
3'h4,
3'h1,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h1,
3'h4,
3'h5,
3'h1,
3'h1,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h1,
3'h4,
3'h4,
3'h4,
3'h1,
3'h4,
3'h4,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h4,
3'h4,
3'h1,
3'h4,
3'h4,
3'h4,
3'h1,
3'h1,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h4,
3'h1,
3'h1,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h1,
3'h4,
3'h4,
3'h1,
3'h1,
3'h4,
3'h4,
3'h1,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h1,
3'h4,
3'h5,
3'h1,
3'h1,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h1,
3'h4,
3'h4,
3'h4,
3'h1,
3'h4,
3'h4,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h4,
3'h4,
3'h1,
3'h4,
3'h4,
3'h4,
3'h1,
3'h1,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h4,
3'h4,
3'h1,
3'h4,
3'h4,
3'h4,
3'h1,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h1,
3'h1,
3'h4,
3'h4,
3'h1,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h1,
3'h1,
3'h4,
3'h1,
3'h1,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h1,
3'h1,
3'h4,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h4,
3'h4,
3'h1,
3'h1,
3'h4,
3'h4,
3'h1,
3'h1,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h4,
3'h1,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h1,
3'h1,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h1,
3'h4,
3'h4,
3'h1,
3'h1,
3'h4,
3'h4,
3'h1,
3'h4,
3'h4,
3'h4,
3'h1,
3'h4,
3'h4,
3'h4,
3'h1,
3'h4,
3'h4,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h4,
3'h4,
3'h1,
3'h4,
3'h4,
3'h4,
3'h1,
3'h1,
3'h4,
3'h4,
3'h1,
3'h4,
3'h1,
3'h1,
3'h4,
3'h1,
3'h1,
3'h4,
3'h4,
3'h1,
3'h4,
3'h4,
3'h4,
3'h1,
3'h4,
3'h4,
3'h4,
3'h1,
3'h4,
3'h4,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h4,
3'h1,
3'h1,
3'h4,
3'h4,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h4,
3'h4,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h4,
3'h4,
3'h4,
3'h1,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h1,
3'h4,
3'h1,
3'h1,
3'h1,
3'h5,
3'h1,
3'h4,
3'h4,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h4,
3'h1,
3'h1,
3'h4,
3'h4,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h4,
3'h4,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h4,
3'h4,
3'h4,
3'h1,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h1,
3'h4,
3'h1,
3'h1,
3'h4,
3'h4,
3'h1,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h1,
3'h1,
3'h4,
3'h1,
3'h1,
3'h1,
3'h4,
3'h1,
3'h1,
3'h4,
3'h4,
3'h4,
3'h1,
3'h4,
3'h4,
3'h1,
3'h1,
3'h4,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h4,
3'h1,
3'h1,
3'h4,
3'h4,
3'h1,
3'h1,
3'h1,
3'h4,
3'h1,
3'h1,
3'h4,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h4,
3'h4,
3'h1,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h1,
3'h4,
3'h1,
3'h1,
3'h1,
3'h4,
3'h4,
3'h1,
3'h4,
3'h4,
3'h4,
3'h1,
3'h1,
3'h1,
3'h1,
3'h4,
3'h1,
3'h1,
3'h1,
3'h4,
3'h1,
3'h4,
3'h4,
3'h4,
3'h1,
3'h4,
3'h4,
3'h4,
3'h1,
3'h4,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h4,
3'h4,
3'h1,
3'h1,
3'h1,
3'h4,
3'h1,
3'h1,
3'h4,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h4,
3'h1,
3'h1,
3'h4,
3'h4,
3'h1,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h1,
3'h4,
3'h4,
3'h1,
3'h1,
3'h4,
3'h4,
3'h1,
3'h1,
3'h4,
3'h4,
3'h4,
3'h1,
3'h1,
3'h1,
3'h4,
3'h1,
3'h1,
3'h4,
3'h4,
3'h1,
3'h4,
3'h4,
3'h4,
3'h1,
3'h4,
3'h4,
3'h4,
3'h1,
3'h4,
3'h4,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h4,
3'h1,
3'h1,
3'h4,
3'h4,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h4,
3'h4,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h4,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h4,
3'h1,
3'h1,
3'h4,
3'h4,
3'h1,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h1,
3'h4,
3'h4,
3'h1,
3'h1,
3'h4,
3'h4,
3'h1,
3'h1,
3'h4,
3'h4,
3'h4,
3'h1,
3'h1,
3'h1,
3'h4,
3'h1,
3'h1,
3'h4,
3'h4,
3'h1,
3'h4,
3'h4,
3'h4,
3'h1,
3'h4,
3'h4,
3'h4,
3'h1,
3'h4,
3'h4,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h4,
3'h1,
3'h1,
3'h4,
3'h4,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h4,
3'h4,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h4,
3'h4,
3'h4,
3'h1,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h1,
3'h4,
3'h1,
3'h1,
3'h4,
3'h4,
3'h1,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h1,
3'h1,
3'h4,
3'h1,
3'h1,
3'h1,
3'h4,
3'h1,
3'h1,
3'h4,
3'h4,
3'h4,
3'h1,
3'h4,
3'h4,
3'h1,
3'h1,
3'h4,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h4,
3'h1,
3'h1,
3'h4,
3'h4,
3'h1,
3'h1,
3'h1,
3'h4,
3'h1,
3'h1,
3'h4,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h4,
3'h4,
3'h1,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h4,
3'h1,
3'h4,
3'h1,
3'h1,
3'h1,
3'h4,
3'h4,
3'h1,
3'h4,
3'h4,
3'h4,
3'h1,
3'h1,
3'h1,
3'h1,
3'h4,
3'h1,
3'h1,
3'h1,
3'h4,
3'h1,
3'h4,
3'h4,
3'h4,
3'h1,
3'h4,
3'h4,
3'h4,
3'h1,
3'h4,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h4,
3'h4,
3'h4,
3'h1,
3'h1,
3'h4,
3'h4,
3'h1,
3'h4,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h4,
3'h4,
3'h1,
3'h1,
3'h4,
3'h4,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h4,
3'h4,
3'h1,
3'h4,
3'h4,
3'h4,
3'h1,
3'h4,
3'h1,
3'h1,
3'h4,
3'h1,
3'h1,
3'h1,
3'h4,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h4,
3'h4,
3'h1,
3'h4,
3'h4,
3'h4,
3'h1,
3'h4,
3'h1,
3'h1,
3'h4,
3'h1,
3'h1,
3'h1,
3'h4,
3'h1,
3'h1,
3'h1,
3'h4,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h4,
3'h4,
3'h4,
3'h1,
3'h4,
3'h4,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h4,
3'h1,
3'h4,
3'h4,
3'h4,
3'h1,
3'h4,
3'h4,
3'h1,
3'h4,
3'h1,
3'h1,
3'h1,
3'h4,
3'h4,
3'h1,
3'h1,
3'h4,
3'h4,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h4,
3'h4,
3'h1,
3'h4,
3'h4,
3'h4,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h4,
3'h1,
3'h1,
3'h4,
3'h4,
3'h1,
3'h4,
3'h4,
3'h1,
3'h4,
3'h4,
3'h1,
3'h1,
3'h4,
3'h4,
3'h1,
3'h1,
3'h4,
3'h4,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h4,
3'h4,
3'h1,
3'h1,
3'h4,
3'h4,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h4,
3'h1,
3'h1,
3'h4,
3'h4,
3'h1,
3'h4,
3'h4,
3'h1,
3'h4,
3'h4,
3'h1,
3'h1,
3'h4,
3'h4,
3'h1,
3'h1,
3'h4,
3'h4,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h4,
3'h4,
3'h1,
3'h1,
3'h4,
3'h4,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h4,
3'h4,
3'h1,
3'h4,
3'h4,
3'h4,
3'h1,
3'h4,
3'h1,
3'h1,
3'h4,
3'h1,
3'h1,
3'h1,
3'h4,
3'h1,
3'h1,
3'h1,
3'h4,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h4,
3'h4,
3'h4,
3'h1,
3'h4,
3'h4,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h4,
3'h1,
3'h4,
3'h4,
3'h4,
3'h1,
3'h4,
3'h4,
3'h1,
3'h4,
3'h1,
3'h1,
3'h1,
3'h4,
3'h4,
3'h1,
3'h1,
3'h4,
3'h4,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h4,
3'h4,
3'h1,
3'h4,
3'h4,
3'h4,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h4,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h4,
3'h1,
3'h1,
3'h4,
3'h4,
3'h1,
3'h4,
3'h1,
3'h1,
3'h4,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h4,
3'h1,
3'h1,
3'h4,
3'h4,
3'h1,
3'h4,
3'h1,
3'h1,
3'h4,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h4,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h4,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h4,
3'h1,
3'h1,
3'h4,
3'h4,
3'h1,
3'h1,
3'h1,
3'h1,
3'h4,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h4,
3'h1,
3'h1,
3'h4,
3'h4,
3'h1,
3'h1,
3'h4,
3'h1,
3'h4,
3'h4,
3'h1,
3'h1,
3'h1,
3'h4,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h4,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h4,
3'h1,
3'h1,
3'h4,
3'h4,
3'h1,
3'h1,
3'h4,
3'h1,
3'h4,
3'h4,
3'h1,
3'h1,
3'h1,
3'h4,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h4,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h4,
3'h1,
3'h1,
3'h4,
3'h4,
3'h1,
3'h4,
3'h1,
3'h1,
3'h4,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h4,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h4,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h4,
3'h1,
3'h1,
3'h4,
3'h4,
3'h1,
3'h1,
3'h1,
3'h1,
3'h4,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h4,
3'h4,
3'h1,
3'h1,
3'h1,
3'h4,
3'h4,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h4,
3'h4,
3'h1,
3'h1,
3'h1,
3'h4,
3'h4,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h4,
3'h1,
3'h1,
3'h1,
3'h4,
3'h1,
3'h1,
3'h1,
3'h1,
3'h4,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h4,
3'h4,
3'h1,
3'h1,
3'h1,
3'h4,
3'h4,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h4,
3'h4,
3'h1,
3'h1,
3'h1,
3'h4,
3'h4,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h4,
3'h4,
3'h1,
3'h1,
3'h1,
3'h4,
3'h4,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h4,
3'h1,
3'h1,
3'h1,
3'h4,
3'h1,
3'h1,
3'h1,
3'h1,
3'h4,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h4,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h4,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1,
3'h1
};

endmodule
