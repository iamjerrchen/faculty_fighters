/* font_rom
 *		This module contains read memory of explicit
 *		enumerations from 0-9, a-z, and A-Z with an extra
 *		bitmap representing a space.
 *
 *		The format of each bitmap:
 *			2 rows top and bottom are empty.
 *			1 column left and right are empty.
 *			Remaining rows and columns represent the bitmap.
 */
module font_rom (	input [9:0] addr,
						output [7:0] data
						);
						
	parameter ADDR_WIDTH = 10; // addressability
	parameter DATA_WIDTH = 8;

	assign data = ROM[addr][7:0];//ROM[addr]; // read bitmap for font
	
	// ROM definition
	parameter [0:2**ADDR_WIDTH-1][DATA_WIDTH-1:0] ROM = {
		// n = x00, 0
		8'b00000000, // 0
		8'b00000000, // 1
		8'b01111110, // 2
		8'b01111110, // 3
		8'b01000010, // 4
		8'b01000010, // 5
		8'b01000010, // 6
		8'b01000010, // 7
		8'b01000010, // 8
		8'b01000010, // 9
		8'b01000010, // a
		8'b01000010, // b
		8'b01111110, // c
		8'b01111110, // d
		8'b00000000, // e
		8'b00000000, // f
		// n = x01, 1
		8'b00000000, // 0
		8'b00000000, // 1
		8'b00011100, // 2
		8'b00111100, // 3
		8'b01101100, // 4
		8'b00001100, // 5
		8'b00001100, // 6
		8'b00001100, // 7
		8'b00001100, // 8
		8'b00001100, // 9
		8'b00001100, // a
		8'b00001100, // b
		8'b01111110, // c
		8'b01111110, // d
		8'b00000000, // e
		8'b00000000, // f
		// n = x02, 2
		8'b00000000, // 0
		8'b00000000, // 1
		8'b00111100, // 2
		8'b01111110, // 3
		8'b01100110, // 4
		8'b01100110, // 5
		8'b00000110, // 6
		8'b00001100, // 7
		8'b00011000, // 8
		8'b00110000, // 9
		8'b01100000, // a
		8'b01100000, // b
		8'b01111110, // c
		8'b01111110, // d
		8'b00000000, // e
		8'b00000000, // f
		// n = x03, 3
		8'b00000000, // 0
		8'b00000000, // 1
		8'b00111100, // 2
		8'b01111110, // 3
		8'b01100110, // 4
		8'b00000110, // 5
		8'b00000110, // 6
		8'b00000110, // 7
		8'b00111100, // 8
		8'b00000110, // 9
		8'b00000110, // a
		8'b01100110, // b
		8'b01111110, // c
		8'b00111100, // d
		8'b00000000, // e
		8'b00000000, // f
		// n = x04, 4
		8'b00000000, // 0
		8'b00000000, // 1
		8'b00000110, // 2
		8'b00001110, // 3
		8'b00011110, // 4
		8'b00110110, // 5
		8'b01100110, // 6
		8'b11000110, // 7
		8'b11111110, // 8
		8'b00000110, // 9
		8'b00000110, // a
		8'b00000110, // b
		8'b00000110, // c
		8'b00000110, // d
		8'b00000000, // e
		8'b00000000, // f
		// n = x05, 5
		8'b00000000, // 0
		8'b00000000, // 1
		8'b01111110, // 2
		8'b01111110, // 3
		8'b01100000, // 4
		8'b01100000, // 5
		8'b01101100, // 6
		8'b01111110, // 7
		8'b01110110, // 8
		8'b00000110, // 9
		8'b00000110, // a
		8'b01100110, // b
		8'b01111110, // c
		8'b00111100, // d
		8'b00000000, // e
		8'b00000000, // f
		// n = x06, 6
		8'b00000000, // 0
		8'b00000000, // 1
		8'b00111100, // 2
		8'b01100110, // 3
		8'b01100110, // 4
		8'b01100110, // 5
		8'b01100000, // 6
		8'b01100000, // 7
		8'b01111000, // 8
		8'b01111110, // 9
		8'b01100110, // a
		8'b01100110, // b
		8'b01100110, // c
		8'b00111100, // d
		8'b00000000, // e
		8'b00000000, // f
		// n = x07, 7
		8'b00000000, // 0
		8'b00000000, // 1
		8'b01111110, // 2
		8'b01111110, // 3
		8'b00000110, // 4
		8'b00001100, // 5
		8'b00011000, // 6
		8'b00011000, // 7
		8'b00110000, // 8
		8'b00110000, // 9
		8'b01100000, // a
		8'b01100000, // b
		8'b01100000, // c
		8'b01100000, // d
		8'b00000000, // e
		8'b00000000, // f
		// n = x08, 8
		8'b00000000, // 0
		8'b00000000, // 1
		8'b00111100, // 2
		8'b01111110, // 3
		8'b01100110, // 4
		8'b01100110, // 5
		8'b01100110, // 6
		8'b00111100, // 7
		8'b00111100, // 8
		8'b01100110, // 9
		8'b01100110, // a
		8'b01100110, // b
		8'b01111110, // c
		8'b00111100, // d
		8'b00000000, // e
		8'b00000000, // f
		// n = x09, 9
		8'b00000000, // 0
		8'b00000000, // 1
		8'b00111100, // 2
		8'b01100110, // 3
		8'b01100110, // 4
		8'b01100110, // 5
		8'b01100110, // 6
		8'b00111110, // 7
		8'b00000110, // 8
		8'b00000110, // 9
		8'b01100110, // a
		8'b01100110, // b
		8'b01100110, // c
		8'b00111110, // d
		8'b00000000, // e
		8'b00000000, // f
		// n = x0A, A
		8'b00000000, // 0
		8'b00000000, // 1
		8'b00011000, // 2
		8'b00111100, // 3
		8'b01111110, // 4
		8'b01100110, // 5
		8'b01100110, // 6
		8'b01100110, // 7
		8'b01111110, // 8
		8'b01111110, // 9
		8'b01100110, // a
		8'b01100110, // b
		8'b01100110, // c
		8'b01100110, // d
		8'b00000000, // e
		8'b00000000, // f
		// n = x0B, B
		8'b00000000, // 0
		8'b00000000, // 1
		8'b01111100, // 2
		8'b01111100, // 3
		8'b01100110, // 4
		8'b01100110, // 5
		8'b01100110, // 6
		8'b01111100, // 7
		8'b01111100, // 8
		8'b01100110, // 9
		8'b01100110, // a
		8'b01100110, // b
		8'b01111100, // c
		8'b01111100, // d
		8'b00000000, // e
		8'b00000000, // f
		// n = x0C, C
		8'b00000000, // 0
		8'b00000000, // 1
		8'b00111100, // 2
		8'b01111110, // 3
		8'b01100110, // 4
		8'b01100110, // 5
		8'b01100000, // 6
		8'b01100000, // 7
		8'b01100000, // 8
		8'b01100000, // 9
		8'b01100110, // a
		8'b01100110, // b
		8'b01111110, // c
		8'b00111100, // d
		8'b00000000, // e
		8'b00000000, // f
		// n = x0D, D
		8'b00000000, // 0
		8'b00000000, // 1
		8'b01111000, // 2
		8'b01111100, // 3
		8'b01100110, // 4
		8'b01100110, // 5
		8'b01100110, // 6
		8'b01100110, // 7
		8'b01100110, // 8
		8'b01100110, // 9
		8'b01100110, // a
		8'b01100110, // b
		8'b01111100, // c
		8'b01111000, // d
		8'b00000000, // e
		8'b00000000, // f
		// n = x0E, E
		8'b00000000, // 0
		8'b00000000, // 1
		8'b01111110, // 2
		8'b01111110, // 3
		8'b01100000, // 4
		8'b01100000, // 5
		8'b01100000, // 6
		8'b01111110, // 7
		8'b01111110, // 8
		8'b01100000, // 9
		8'b01100000, // a
		8'b01100000, // b
		8'b01111110, // c
		8'b01111110, // d
		8'b00000000, // e
		8'b00000000, // f
		// n = x0F, F
		8'b00000000, // 0
		8'b00000000, // 1
		8'b01111110, // 2
		8'b01111110, // 3
		8'b01100000, // 4
		8'b01100000, // 5
		8'b01100000, // 6
		8'b01111110, // 7
		8'b01111110, // 8
		8'b01100000, // 9
		8'b01100000, // a
		8'b01100000, // b
		8'b01100000, // c
		8'b01100000, // d
		8'b00000000, // e
		8'b00000000, // f
		// n = x10, G
		8'b00000000, // 0
		8'b00000000, // 1
		8'b00111100, // 2
		8'b01111110, // 3
		8'b01100110, // 4
		8'b01100000, // 5
		8'b01100000, // 6
		8'b01100000, // 7
		8'b01101110, // 8
		8'b01101110, // 9
		8'b01100110, // a
		8'b01100110, // b
		8'b01111110, // c
		8'b00111110, // d
		8'b00000000, // e
		8'b00000000, // f
		// n = x11, H
		8'b00000000, // 0
		8'b00000000, // 1
		8'b01100110, // 2
		8'b01100110, // 3
		8'b01100110, // 4
		8'b01100110, // 5
		8'b01100110, // 6
		8'b01111110, // 7
		8'b01111110, // 8
		8'b01100110, // 9
		8'b01100110, // a
		8'b01100110, // b
		8'b01100110, // c
		8'b01100110, // d
		8'b00000000, // e
		8'b00000000, // f
		// n = x12, I
		8'b00000000, // 0
		8'b00000000, // 1
		8'b01111110, // 2
		8'b01111110, // 3
		8'b00011000, // 4
		8'b00011000, // 5
		8'b00011000, // 6
		8'b00011000, // 7
		8'b00011000, // 8
		8'b00011000, // 9
		8'b00011000, // a
		8'b00011000, // b
		8'b01111110, // c
		8'b01111110, // d
		8'b00000000, // e
		8'b00000000, // f
		// n = x13, J
		8'b00000000, // 0
		8'b00000000, // 1
		8'b01111111, // 2
		8'b01111111, // 3
		8'b00001100, // 4
		8'b00001100, // 5
		8'b00001100, // 6
		8'b00001100, // 7
		8'b00001100, // 8
		8'b01101100, // 9
		8'b01101100, // a
		8'b01101100, // b
		8'b01111100, // c
		8'b00111000, // d
		8'b00000000, // e
		8'b00000000, // f
		// n = x14, K
		8'b00000000, // 0
		8'b00000000, // 1
		8'b01100110, // 2
		8'b01100110, // 3
		8'b01100110, // 4
		8'b01101100, // 5
		8'b01101100, // 6
		8'b01111000, // 7
		8'b01111000, // 8
		8'b01101100, // 9
		8'b01101100, // a
		8'b01100110, // b
		8'b01100110, // c
		8'b01100110, // d
		8'b00000000, // e
		8'b00000000, // f
		// n = x15, L
		8'b00000000, // 0
		8'b00000000, // 1
		8'b01100000, // 2
		8'b01100000, // 3
		8'b01100000, // 4
		8'b01100000, // 5
		8'b01100000, // 6
		8'b01100000, // 7
		8'b01100000, // 8
		8'b01100000, // 9
		8'b01100000, // a
		8'b01100000, // b
		8'b01111110, // c
		8'b01111110, // d
		8'b00000000, // e
		8'b00000000, // f
		// n = x16, M
		8'b00000000, // 0
		8'b00000000, // 1
		8'b01000010, // 2
		8'b01000010, // 3
		8'b01100110, // 4
		8'b01100110, // 5
		8'b01111110, // 6
		8'b01011010, // 7
		8'b01011010, // 8
		8'b01000010, // 9
		8'b01000010, // a
		8'b01000010, // b
		8'b01000010, // c
		8'b01000010, // d
		8'b00000000, // e
		8'b00000000, // f
		// n = x17, N
		8'b00000000, // 0
		8'b00000000, // 1
		8'b01100110, // 2
		8'b01100110, // 3
		8'b01100110, // 4
		8'b01110110, // 5
		8'b01110110, // 6
		8'b01111110, // 7
		8'b01111110, // 8
		8'b01101110, // 9
		8'b01101110, // a
		8'b01100110, // b
		8'b01100110, // c
		8'b01100110, // d
		8'b00000000, // e
		8'b00000000, // f
		// n = x18, O
		8'b00000000, // 0
		8'b00000000, // 1
		8'b00111100, // 2
		8'b01111110, // 3
		8'b01100110, // 4
		8'b01100110, // 5
		8'b01100110, // 6
		8'b01100110, // 7
		8'b01100110, // 8
		8'b01100110, // 9
		8'b01100110, // a
		8'b01100110, // b
		8'b01111110, // c
		8'b00111100, // d
		8'b00000000, // e
		8'b00000000, // f
		// n = x19, P
		8'b00000000, // 0
		8'b00000000, // 1
		8'b0111110, // 2
		8'b01111110, // 3
		8'b01100110, // 4
		8'b01100110, // 5
		8'b01100110, // 6
		8'b01111110, // 7
		8'b01111100, // 8
		8'b01100000, // 9
		8'b01100000, // a
		8'b01100000, // b
		8'b01100000, // c
		8'b01100000, // d
		8'b00000000, // e
		8'b00000000, // f
		// n = x1A, Q
		8'b00000000, // 0
		8'b00000000, // 1
		8'b00111000, // 2
		8'b01111100, // 3
		8'b01100100, // 4
		8'b01100100, // 5
		8'b01100100, // 6
		8'b01100100, // 7
		8'b01100100, // 8
		8'b01100100, // 9
		8'b01100100, // a
		8'b01100100, // b
		8'b01100100, // c
		8'b00111110, // d
		8'b00000000, // e
		8'b00000000, // f
		// n = x1B, R
		8'b00000000, // 0
		8'b00000000, // 1
		8'b01111100, // 2
		8'b01111110, // 3
		8'b01100110, // 4
		8'b01100110, // 5
		8'b01100110, // 6
		8'b01111110, // 7
		8'b01111100, // 8
		8'b01101100, // 9
		8'b01101100, // a
		8'b01100110, // b
		8'b01100110, // c
		8'b01100110, // d
		8'b00000000, // e
		8'b00000000, // f
		// n = x1C, S
		8'b00000000, // 0
		8'b00000000, // 1
		8'b00111100, // 2
		8'b01111110, // 3
		8'b01100110, // 4
		8'b01100010, // 5
		8'b01100000, // 6
		8'b01111100, // 7
		8'b00111110, // 8
		8'b00000110, // 9
		8'b01000110, // a
		8'b01100110, // b
		8'b01111110, // c
		8'b00111100, // d
		8'b00000000, // e
		8'b00000000, // f
		// n = x1D, T
		8'b00000000, // 0
		8'b00000000, // 1
		8'b01111110, // 2
		8'b01111110, // 3
		8'b00011000, // 4
		8'b00011000, // 5
		8'b00011000, // 6
		8'b00011000, // 7
		8'b00011000, // 8
		8'b00011000, // 9
		8'b00011000, // a
		8'b00011000, // b
		8'b00011000, // c
		8'b00011000, // d
		8'b00000000, // e
		8'b00000000, // f
		// n = x1E, U
		8'b00000000, // 0
		8'b00000000, // 1
		8'b01100110, // 2
		8'b01100110, // 3
		8'b01100110, // 4
		8'b01100110, // 5
		8'b01100110, // 6
		8'b01100110, // 7
		8'b01100110, // 8
		8'b01100110, // 9
		8'b01100110, // a
		8'b01100110, // b
		8'b01111110, // c
		8'b00111100, // d
		8'b00000000, // e
		8'b00000000, // f
		// n = x1F, V
		8'b00000000, // 0
		8'b00000000, // 1
		8'b01100110, // 2
		8'b01100110, // 3
		8'b01100110, // 4
		8'b01100110, // 5
		8'b01100110, // 6
		8'b01100110, // 7
		8'b01100110, // 8
		8'b01100110, // 9
		8'b01111110, // a
		8'b00111100, // b
		8'b00011000, // c
		8'b00011000, // d
		8'b00000000, // e
		8'b00000000, // f
		// n = x20, W
		8'b00000000, // 0
		8'b00000000, // 1
		8'b01000010, // 2
		8'b01000010, // 3
		8'b01000010, // 4
		8'b01000010, // 5
		8'b01000010, // 6
		8'b01000010, // 7
		8'b01011010, // 8
		8'b01011010, // 9
		8'b01111110, // a
		8'b01100110, // b
		8'b01100110, // c
		8'b01000010, // d
		8'b00000000, // e
		8'b00000000, // f
		// n = x21, X
		8'b00000000, // 0
		8'b00000000, // 1
		8'b01100110, // 2
		8'b01100110, // 3
		8'b01100110, // 4
		8'b01100110, // 5
		8'b00111100, // 6
		8'b00011000, // 7
		8'b00011000, // 8
		8'b00111100, // 9
		8'b01100110, // a
		8'b01100110, // b
		8'b01100110, // c
		8'b01100110, // d
		8'b00000000, // e
		8'b00000000, // f
		// n = x22, Y
		8'b00000000, // 0
		8'b00000000, // 1
		8'b01100110, // 2
		8'b01100110, // 3
		8'b01100110, // 4
		8'b01100110, // 5
		8'b00111100, // 6
		8'b00111100, // 7
		8'b00011000, // 8
		8'b00011000, // 9
		8'b00011000, // a
		8'b00011000, // b
		8'b00011000, // c
		8'b00011000, // d
		8'b00000000, // e
		8'b00000000, // f
		// n = x23, Z
		8'b00000000, // 0
		8'b00000000, // 1
		8'b01111110, // 2
		8'b01111110, // 3
		8'b00000110, // 4
		8'b00000110, // 5
		8'b00001100, // 6
		8'b00001100, // 7
		8'b00011000, // 8
		8'b00110000, // 9
		8'b00110000, // a
		8'b01100000, // b
		8'b01111110, // c
		8'b01111110, // d
		8'b00000000, // e
		8'b00000000, // f
		// n = x24, a
		8'b00000000, // 0
		8'b00000000, // 1
		8'b00000000, // 2
		8'b00000000, // 3
		8'b00000000, // 4
		8'b00000000, // 5
		8'b00000000, // 6
		8'b00000000, // 7
		8'b00111000, // 8
		8'b01101100, // 9
		8'b01101100, // a
		8'b01101110, // b
		8'b01101110, // c
		8'b00111010, // d
		8'b00000000, // e
		8'b00000000, // f
		// n = x25, b
		8'b00000000, // 0
		8'b00000000, // 1
		8'b00000000, // 2
		8'b01100000, // 3
		8'b01100000, // 4
		8'b01100000, // 5
		8'b01100000, // 6
		8'b01100000, // 7
		8'b01111100, // 8
		8'b01100110, // 9
		8'b01100110, // a
		8'b01100110, // b
		8'b01100110, // c
		8'b01111100, // d
		8'b00000000, // e
		8'b00000000, // f
		// n = x26, c
		8'b00000000, // 0
		8'b00000000, // 1
		8'b00000000, // 2
		8'b00000000, // 3
		8'b00000000, // 4
		8'b00000000, // 5
		8'b00000000, // 6
		8'b00000000, // 7
		8'b00111100, // 8
		8'b01100110, // 9
		8'b01100000, // a
		8'b01100000, // b
		8'b01100110, // c
		8'b00111100, // d
		8'b00000000, // e
		8'b00000000, // f
		// n = x27, d
		8'b00000000, // 0
		8'b00000000, // 1
		8'b00000000, // 2
		8'b00000110, // 3
		8'b00000110, // 4
		8'b00000110, // 5
		8'b00000110, // 6
		8'b00000110, // 7
		8'b00111110, // 8
		8'b01100110, // 9
		8'b01100110, // a
		8'b01100110, // b
		8'b01100110, // c
		8'b00111110, // d
		8'b00000000, // e
		8'b00000000, // f
		// n = x28, e
		8'b00000000, // 0
		8'b00000000, // 1
		8'b00000000, // 2
		8'b00000000, // 3
		8'b00000000, // 4
		8'b00000000, // 5
		8'b00000000, // 6
		8'b00000000, // 7
		8'b00111100, // 8
		8'b01100110, // 9
		8'b01111110, // a
		8'b01100000, // b
		8'b01100000, // c
		8'b00111100, // d
		8'b00000000, // e
		8'b00000000, // f
		// n = x29, f
		8'b00000000, // 0
		8'b00000000, // 1
		8'b00000000, // 2
		8'b00011100, // 3
		8'b00111110, // 4
		8'b00110110, // 5
		8'b00110110, // 6
		8'b00110000, // 7
		8'b00110000, // 8
		8'b01111100, // 9
		8'b01111100, // a
		8'b00110000, // b
		8'b00110000, // c
		8'b00110000, // d
		8'b00000000, // e
		8'b00000000, // f
		// n = x2A, g
		8'b00000000, // 0
		8'b00000000, // 1
		8'b00000000, // 2
		8'b00000000, // 3
		8'b00000000, // 4
		8'b00000000, // 5
		8'b00000000, // 6
		8'b00000000, // 7
		8'b00111100, // 8
		8'b01100110, // 9
		8'b01100110, // a
		8'b01111110, // b
		8'b00000110, // c
		8'b00000110, // d
		8'b00000110, // e
		8'b01111100, // f
		// n = x2B, h
		8'b00000000, // 0
		8'b00000000, // 1
		8'b00000000, // 2
		8'b01100000, // 3
		8'b01100000, // 4
		8'b01100000, // 5
		8'b01100000, // 6
		8'b01100000, // 7
		8'b01101100, // 8
		8'b01111110, // 9
		8'b01100110, // a
		8'b01100110, // b
		8'b01100110, // c
		8'b01100110, // d
		8'b00000000, // e
		8'b00000000, // f
		// n = x2C, i
		8'b00000000, // 0
		8'b00000000, // 1
		8'b00000000, // 2
		8'b00011000, // 3
		8'b00111100, // 4
		8'b00111100, // 5
		8'b00011000, // 6
		8'b00000000, // 7
		8'b00011000, // 8
		8'b00011000, // 9
		8'b00011000, // a
		8'b00011000, // b
		8'b00011000, // c
		8'b00011000, // d
		8'b00000000, // e
		8'b00000000, // f
		// n = x2D, j
		8'b00000000, // 0
		8'b00000000, // 1
		8'b00000000, // 2
		8'b00001100, // 3
		8'b00011110, // 4
		8'b00011110, // 5
		8'b00001100, // 6
		8'b00000000, // 7
		8'b00001100, // 8
		8'b00001100, // 9
		8'b00001100, // a
		8'b00001100, // b
		8'b01101100, // c
		8'b01101100, // d
		8'b01101100, // e
		8'b01111100, // f
		// n = x2E, k
		8'b00000000, // 0
		8'b00000000, // 1
		8'b00000000, // 2
		8'b01100000, // 3
		8'b01100000, // 4
		8'b01100000, // 5
		8'b01100000, // 6
		8'b01100000, // 7
		8'b01100110, // 8
		8'b01101100, // 9
		8'b01111000, // a
		8'b01111000, // b
		8'b01101100, // c
		8'b01100110, // d
		8'b00000000, // e
		8'b00000000, // f
		// n = x2F, l
		8'b00000000, // 0
		8'b00000000, // 1
		8'b00000000, // 2
		8'b00011000, // 3
		8'b00011000, // 4
		8'b00011000, // 5
		8'b00011000, // 6
		8'b00011000, // 7
		8'b00011000, // 8
		8'b00011000, // 9
		8'b00011000, // a
		8'b00011000, // b
		8'b00011000, // c
		8'b00011000, // d
		8'b00000000, // e
		8'b00000000, // f
		// n = x30, m
		8'b00000000, // 0
		8'b00000000, // 1
		8'b00000000, // 2
		8'b00000000, // 3
		8'b00000000, // 4
		8'b00000000, // 5
		8'b00000000, // 6
		8'b00000000, // 7
		8'b00100100, // 8
		8'b01011010, // 9
		8'b01011010, // a
		8'b01011010, // b
		8'b01011010, // c
		8'b01000010, // d
		8'b00000000, // e
		8'b00000000, // f
		// n = x31, n
		8'b00000000, // 0
		8'b00000000, // 1
		8'b00000000, // 2
		8'b00000000, // 3
		8'b00000000, // 4
		8'b00000000, // 5
		8'b00000000, // 6
		8'b00000000, // 7
		8'b00011000, // 8
		8'b00111100, // 9
		8'b01100110, // a
		8'b01100110, // b
		8'b01100110, // c
		8'b01100110, // d
		8'b00000000, // e
		8'b00000000, // f
		// n = x32, o
		8'b00000000, // 0
		8'b00000000, // 1
		8'b00000000, // 2
		8'b00000000, // 3
		8'b00000000, // 4
		8'b00000000, // 5
		8'b00000000, // 6
		8'b00000000, // 7
		8'b00111100, // 8
		8'b01111110, // 9
		8'b01100110, // a
		8'b01100110, // b
		8'b01111110, // c
		8'b00111100, // d
		8'b00000000, // e
		8'b00000000, // f
		// n = x33, p
		8'b00000000, // 0
		8'b00000000, // 1
		8'b00000000, // 2
		8'b00000000, // 3
		8'b00000000, // 4
		8'b00000000, // 5
		8'b00000000, // 6
		8'b00000000, // 7
		8'b00111100, // 8
		8'b01100110, // 9
		8'b01100110, // a
		8'b01100110, // b
		8'b01111100, // c
		8'b01100000, // d
		8'b01100000, // e
		8'b01100000, // f
		// n = x34, q
		8'b00000000, // 0
		8'b00000000, // 1
		8'b00000000, // 2
		8'b00000000, // 3
		8'b00000000, // 4
		8'b00000000, // 5
		8'b00000000, // 6
		8'b00000000, // 7
		8'b00111100, // 8
		8'b01100110, // 9
		8'b01100110, // a
		8'b01100110, // b
		8'b00111110, // c
		8'b00000110, // d
		8'b00000110, // e
		8'b00000110, // f
		// n = x35, r
		8'b00000000, // 0
		8'b00000000, // 1
		8'b00000000, // 2
		8'b00000000, // 3
		8'b00000000, // 4
		8'b00000000, // 5
		8'b00000000, // 6
		8'b00000000, // 7
		8'b01001110, // 8
		8'b01111000, // 9
		8'b01100000, // a
		8'b01000000, // b
		8'b01000000, // c
		8'b01000000, // d
		8'b00000000, // e
		8'b00000000, // f
		// n = x36, s
		8'b00000000, // 0
		8'b00000000, // 1
		8'b00000000, // 2
		8'b00000000, // 3
		8'b00000000, // 4
		8'b00000000, // 5
		8'b00000000, // 6
		8'b00111100, // 7
		8'b01100110, // 8
		8'b01100000, // 9
		8'b00111100, // a
		8'b00000110, // b
		8'b01100110, // c
		8'b00111100, // d
		8'b00000000, // e
		8'b00000000, // f
		// n = x37, t
		8'b00000000, // 0
		8'b00000000, // 1
		8'b00000000, // 2
		8'b00011000, // 3
		8'b00011000, // 4
		8'b00011000, // 5
		8'b00011000, // 6
		8'b01111110, // 7
		8'b01111110, // 8
		8'b00011000, // 9
		8'b00011000, // a
		8'b00011000, // b
		8'b00011000, // c
		8'b00011000, // d
		8'b00000000, // e
		8'b00000000, // f
		// n = x38, u
		8'b00000000, // 0
		8'b00000000, // 1
		8'b00000000, // 2
		8'b00000000, // 3
		8'b00000000, // 4
		8'b00000000, // 5
		8'b00000000, // 6
		8'b01100110, // 7
		8'b01100110, // 8
		8'b01100110, // 9
		8'b01100110, // a
		8'b01100110, // b
		8'b01111110, // c
		8'b00111010, // d
		8'b00000000, // e
		8'b00000000, // f
		// n = x39, v
		8'b00000000, // 0
		8'b00000000, // 1
		8'b00000000, // 2
		8'b00000000, // 3
		8'b00000000, // 4
		8'b00000000, // 5
		8'b00000000, // 6
		8'b00000000, // 7
		8'b01100110, // 8
		8'b01100110, // 9
		8'b01100110, // a
		8'b01100110, // b
		8'b00111100, // c
		8'b00011000, // d
		8'b00000000, // e
		8'b00000000, // f
		// n = x3A, w
		8'b00000000, // 0
		8'b00000000, // 1
		8'b00000000, // 2
		8'b00000000, // 3
		8'b00000000, // 4
		8'b00000000, // 5
		8'b00000000, // 6
		8'b00000000, // 7
		8'b01000010, // 8
		8'b01000010, // 9
		8'b01011010, // a
		8'b01011010, // b
		8'b01011010, // c
		8'b00100100, // d
		8'b00000000, // e
		8'b00000000, // f
		// n = x3B, x
		8'b00000000, // 0
		8'b00000000, // 1
		8'b00000000, // 2
		8'b00000000, // 3
		8'b00000000, // 4
		8'b00000000, // 5
		8'b00000000, // 6
		8'b00000000, // 7
		8'b01100110, // 8
		8'b01100110, // 9
		8'b00111100, // a
		8'b00111100, // b
		8'b01100110, // c
		8'b01100110, // d
		8'b00000000, // e
		8'b00000000, // f
		// n = x3C, y
		8'b00000000, // 0
		8'b00000000, // 1
		8'b00000000, // 2
		8'b00000000, // 3
		8'b00000000, // 4
		8'b00000000, // 5
		8'b00000000, // 6
		8'b00000000, // 7
		8'b01100110, // 8
		8'b01100110, // 9
		8'b01100110, // a
		8'b01100110, // b
		8'b01111110, // c
		8'b00000110, // d
		8'b00000110, // e
		8'b00000110, // f
		// n = x3D, z
		8'b00000000, // 0
		8'b00000000, // 1
		8'b00000000, // 2
		8'b00000000, // 3
		8'b00000000, // 4
		8'b00000000, // 5
		8'b00000000, // 6
		8'b01111110, // 7
		8'b00000110, // 8
		8'b00001100, // 9
		8'b00011000, // a
		8'b00110000, // b
		8'b01100000, // c
		8'b01111110, // d
		8'b00000000, // e
		8'b00000000, // f
		// n = x3E, space
		8'b00000000, // 0
		8'b00000000, // 1
		8'b00000000, // 2
		8'b00000000, // 3
		8'b00000000, // 4
		8'b00000000, // 5
		8'b00000000, // 6
		8'b00000000, // 7
		8'b00000000, // 8
		8'b00000000, // 9
		8'b00000000, // a
		8'b00000000, // b
		8'b00000000, // c
		8'b00000000, // d
		8'b00000000, // e
		8'b00000000, // f
		// n = x3F, !
		8'b00000000, // 0
		8'b00110000, // 1
		8'b01111000, // 2
		8'b01111000, // 3
		8'b01111000, // 4
		8'b01111000, // 5
		8'b01111000, // 6
		8'b01111000, // 7
		8'b01111000, // 8
		8'b01111000, // 9
		8'b00110000, // a
		8'b00000000, // b
		8'b00110000, // c
		8'b00110000, // d
		8'b00000000, // e
		8'b00000000  // f
	};

			
endmodule
